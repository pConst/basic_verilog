
`ifndef TITLE
`define TITLE "title"
`endif

module one;

initial $display(`TITLE);

endmodule
