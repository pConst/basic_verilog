// Copyright 2007 Altera Corporation. All rights reserved.  
// Altera products are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.  
//
// This reference design file, and your use thereof, is subject to and governed
// by the terms and conditions of the applicable Altera Reference Design 
// License Agreement (either as signed by you or found at www.altera.com).  By
// using this reference design file, you indicate your acceptance of such terms
// and conditions between you and Altera Corporation.  In the event that you do
// not agree with such terms and conditions, you may not use the reference 
// design file and please promptly destroy any copies you have made.
//
// This reference design file is being provided on an "as-is" basis and as an 
// accommodation and therefore all warranties, representations or guarantees of 
// any kind (whether express, implied or statutory) including, without 
// limitation, warranties of merchantability, non-infringement, or fitness for
// a particular purpose, are specifically disclaimed.  By making this reference
// design file available, Altera expressly does not recommend, suggest or 
// require that this reference design file be used in combination with any 
// other product not provided by Altera.
/////////////////////////////////////////////////////////////////////////////

module mask_32 (in,mask);
input [4:0] in;
output [31:0] mask;
reg [31:0] mask;

parameter FROM_MSB = 1'b1;
parameter DIAG_ONES = 1'b1;

generate
  if (!FROM_MSB && !DIAG_ONES) begin
    always @(in) begin
    case (in)
      5'd0: mask=32'b00000000000000000000000000000000;
      5'd1: mask=32'b00000000000000000000000000000001;
      5'd2: mask=32'b00000000000000000000000000000011;
      5'd3: mask=32'b00000000000000000000000000000111;
      5'd4: mask=32'b00000000000000000000000000001111;
      5'd5: mask=32'b00000000000000000000000000011111;
      5'd6: mask=32'b00000000000000000000000000111111;
      5'd7: mask=32'b00000000000000000000000001111111;
      5'd8: mask=32'b00000000000000000000000011111111;
      5'd9: mask=32'b00000000000000000000000111111111;
      5'd10: mask=32'b00000000000000000000001111111111;
      5'd11: mask=32'b00000000000000000000011111111111;
      5'd12: mask=32'b00000000000000000000111111111111;
      5'd13: mask=32'b00000000000000000001111111111111;
      5'd14: mask=32'b00000000000000000011111111111111;
      5'd15: mask=32'b00000000000000000111111111111111;
      5'd16: mask=32'b00000000000000001111111111111111;
      5'd17: mask=32'b00000000000000011111111111111111;
      5'd18: mask=32'b00000000000000111111111111111111;
      5'd19: mask=32'b00000000000001111111111111111111;
      5'd20: mask=32'b00000000000011111111111111111111;
      5'd21: mask=32'b00000000000111111111111111111111;
      5'd22: mask=32'b00000000001111111111111111111111;
      5'd23: mask=32'b00000000011111111111111111111111;
      5'd24: mask=32'b00000000111111111111111111111111;
      5'd25: mask=32'b00000001111111111111111111111111;
      5'd26: mask=32'b00000011111111111111111111111111;
      5'd27: mask=32'b00000111111111111111111111111111;
      5'd28: mask=32'b00001111111111111111111111111111;
      5'd29: mask=32'b00011111111111111111111111111111;
      5'd30: mask=32'b00111111111111111111111111111111;
      5'd31: mask=32'b01111111111111111111111111111111;
      default: mask=0;
    endcase
    end
  end
  else if ( FROM_MSB && !DIAG_ONES) begin
    always @(in) begin
    case (in)
      5'd0: mask=32'b00000000000000000000000000000000;
      5'd1: mask=32'b10000000000000000000000000000000;
      5'd2: mask=32'b11000000000000000000000000000000;
      5'd3: mask=32'b11100000000000000000000000000000;
      5'd4: mask=32'b11110000000000000000000000000000;
      5'd5: mask=32'b11111000000000000000000000000000;
      5'd6: mask=32'b11111100000000000000000000000000;
      5'd7: mask=32'b11111110000000000000000000000000;
      5'd8: mask=32'b11111111000000000000000000000000;
      5'd9: mask=32'b11111111100000000000000000000000;
      5'd10: mask=32'b11111111110000000000000000000000;
      5'd11: mask=32'b11111111111000000000000000000000;
      5'd12: mask=32'b11111111111100000000000000000000;
      5'd13: mask=32'b11111111111110000000000000000000;
      5'd14: mask=32'b11111111111111000000000000000000;
      5'd15: mask=32'b11111111111111100000000000000000;
      5'd16: mask=32'b11111111111111110000000000000000;
      5'd17: mask=32'b11111111111111111000000000000000;
      5'd18: mask=32'b11111111111111111100000000000000;
      5'd19: mask=32'b11111111111111111110000000000000;
      5'd20: mask=32'b11111111111111111111000000000000;
      5'd21: mask=32'b11111111111111111111100000000000;
      5'd22: mask=32'b11111111111111111111110000000000;
      5'd23: mask=32'b11111111111111111111111000000000;
      5'd24: mask=32'b11111111111111111111111100000000;
      5'd25: mask=32'b11111111111111111111111110000000;
      5'd26: mask=32'b11111111111111111111111111000000;
      5'd27: mask=32'b11111111111111111111111111100000;
      5'd28: mask=32'b11111111111111111111111111110000;
      5'd29: mask=32'b11111111111111111111111111111000;
      5'd30: mask=32'b11111111111111111111111111111100;
      5'd31: mask=32'b11111111111111111111111111111110;
      default: mask=0;
    endcase
    end
  end
  else if (!FROM_MSB &&  DIAG_ONES) begin
    always @(in) begin
    case (in)
      5'd0: mask=32'b00000000000000000000000000000001;
      5'd1: mask=32'b00000000000000000000000000000011;
      5'd2: mask=32'b00000000000000000000000000000111;
      5'd3: mask=32'b00000000000000000000000000001111;
      5'd4: mask=32'b00000000000000000000000000011111;
      5'd5: mask=32'b00000000000000000000000000111111;
      5'd6: mask=32'b00000000000000000000000001111111;
      5'd7: mask=32'b00000000000000000000000011111111;
      5'd8: mask=32'b00000000000000000000000111111111;
      5'd9: mask=32'b00000000000000000000001111111111;
      5'd10: mask=32'b00000000000000000000011111111111;
      5'd11: mask=32'b00000000000000000000111111111111;
      5'd12: mask=32'b00000000000000000001111111111111;
      5'd13: mask=32'b00000000000000000011111111111111;
      5'd14: mask=32'b00000000000000000111111111111111;
      5'd15: mask=32'b00000000000000001111111111111111;
      5'd16: mask=32'b00000000000000011111111111111111;
      5'd17: mask=32'b00000000000000111111111111111111;
      5'd18: mask=32'b00000000000001111111111111111111;
      5'd19: mask=32'b00000000000011111111111111111111;
      5'd20: mask=32'b00000000000111111111111111111111;
      5'd21: mask=32'b00000000001111111111111111111111;
      5'd22: mask=32'b00000000011111111111111111111111;
      5'd23: mask=32'b00000000111111111111111111111111;
      5'd24: mask=32'b00000001111111111111111111111111;
      5'd25: mask=32'b00000011111111111111111111111111;
      5'd26: mask=32'b00000111111111111111111111111111;
      5'd27: mask=32'b00001111111111111111111111111111;
      5'd28: mask=32'b00011111111111111111111111111111;
      5'd29: mask=32'b00111111111111111111111111111111;
      5'd30: mask=32'b01111111111111111111111111111111;
      5'd31: mask=32'b11111111111111111111111111111111;
      default: mask=0;
    endcase
    end
  end
  else if ( FROM_MSB &&  DIAG_ONES) begin
    always @(in) begin
    case (in)
      5'd0: mask=32'b10000000000000000000000000000000;
      5'd1: mask=32'b11000000000000000000000000000000;
      5'd2: mask=32'b11100000000000000000000000000000;
      5'd3: mask=32'b11110000000000000000000000000000;
      5'd4: mask=32'b11111000000000000000000000000000;
      5'd5: mask=32'b11111100000000000000000000000000;
      5'd6: mask=32'b11111110000000000000000000000000;
      5'd7: mask=32'b11111111000000000000000000000000;
      5'd8: mask=32'b11111111100000000000000000000000;
      5'd9: mask=32'b11111111110000000000000000000000;
      5'd10: mask=32'b11111111111000000000000000000000;
      5'd11: mask=32'b11111111111100000000000000000000;
      5'd12: mask=32'b11111111111110000000000000000000;
      5'd13: mask=32'b11111111111111000000000000000000;
      5'd14: mask=32'b11111111111111100000000000000000;
      5'd15: mask=32'b11111111111111110000000000000000;
      5'd16: mask=32'b11111111111111111000000000000000;
      5'd17: mask=32'b11111111111111111100000000000000;
      5'd18: mask=32'b11111111111111111110000000000000;
      5'd19: mask=32'b11111111111111111111000000000000;
      5'd20: mask=32'b11111111111111111111100000000000;
      5'd21: mask=32'b11111111111111111111110000000000;
      5'd22: mask=32'b11111111111111111111111000000000;
      5'd23: mask=32'b11111111111111111111111100000000;
      5'd24: mask=32'b11111111111111111111111110000000;
      5'd25: mask=32'b11111111111111111111111111000000;
      5'd26: mask=32'b11111111111111111111111111100000;
      5'd27: mask=32'b11111111111111111111111111110000;
      5'd28: mask=32'b11111111111111111111111111111000;
      5'd29: mask=32'b11111111111111111111111111111100;
      5'd30: mask=32'b11111111111111111111111111111110;
      5'd31: mask=32'b11111111111111111111111111111111;
      default: mask=0;
    endcase
    end
  end
endgenerate
endmodule
