//------------------------------------------------------------------------------
// fifo_single_clock_reg_v1_init.svh
// published as part of https://github.com/pConst/basic_verilog
// Konstantin Pavlov, pavlovconst@gmail.com
//------------------------------------------------------------------------------

// INFO ------------------------------------------------------------------------
//  Initialization statements example for fifo_single_clock_reg_v1 fifo
//

  data[0] <=  32'hAAAA;
  data[1] <=  32'h0001;
  data[2] <=  32'h0002;
  data[3] <=  32'h0003;
  data[4] <=  32'h0004;
  data[5] <=  32'h0005;
  data[6] <=  32'h0006;
  data[7] <=  32'h0007;
  data[8] <=  32'hBBBB;
  data[9] <=  32'h0001;
  data[10] <= 32'h0002;
  data[11] <= 32'h0003;
  data[12] <= 32'h0004;
  data[13] <= 32'h0005;
  data[14] <= 32'h0006;
  data[15] <= 32'h0007;
  data[16] <= 32'hCCCC;
  data[17] <= 32'h0001;
  data[18] <= 32'h0002;
  data[19] <= 32'h0003;
  data[20] <= 32'h0004;
  data[21] <= 32'h0005;
  data[22] <= 32'h0006;
  data[23] <= 32'h0007;
  data[24] <= 32'hDDDD;
  data[25] <= 32'h0001;
  data[26] <= 32'h0002;
  data[27] <= 32'h0003;
  data[28] <= 32'h0004;
  data[29] <= 32'h0005;
  data[30] <= 32'h0006;
  data[31] <= 32'h0007;

