// Copyright 2007 Altera Corporation. All rights reserved.  
// Altera products are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.  
//
// This reference design file, and your use thereof, is subject to and governed
// by the terms and conditions of the applicable Altera Reference Design 
// License Agreement (either as signed by you or found at www.altera.com).  By
// using this reference design file, you indicate your acceptance of such terms
// and conditions between you and Altera Corporation.  In the event that you do
// not agree with such terms and conditions, you may not use the reference 
// design file and please promptly destroy any copies you have made.
//
// This reference design file is being provided on an "as-is" basis and as an 
// accommodation and therefore all warranties, representations or guarantees of 
// any kind (whether express, implied or statutory) including, without 
// limitation, warranties of merchantability, non-infringement, or fitness for
// a particular purpose, are specifically disclaimed.  By making this reference
// design file available, Altera expressly does not recommend, suggest or 
// require that this reference design file be used in combination with any 
// other product not provided by Altera.
/////////////////////////////////////////////////////////////////////////////

// baeckler - 02-14-2007

module rgb_to_hue (
	clk,rst,
	r,g,b,
	hue
);

input clk,rst;
input [7:0] r,g,b;
output [7:0] hue;

reg [7:0] hue;

wire r_ge_b = (r >= b);
wire r_ge_g = (r >= g);
wire g_ge_b = (g >= b);
wire g_ge_r = (g >= r);
wire b_ge_r = (b >= r);
wire b_ge_g = (b >= g);

reg [7:0] diff_a,diff_b;
reg [3:0] hue_ofs;
reg sub;

always @(posedge clk) begin
	sub <= 1'b0;
	if (r_ge_b & r_ge_g & g_ge_b) begin
		// R G B
		hue_ofs <= 4'h0;
		diff_a <= g - b;
		diff_b <= r - b;
	end
	else if (b_ge_r & g_ge_b & g_ge_r) begin
		// G B R
		hue_ofs <= 4'h5;
		diff_a <= b - r;
		diff_b <= g - r;
	end
	else if (r_ge_b & g_ge_r & g_ge_b) begin
		// G R B
		hue_ofs <= 4'h5;
		sub <= 1'b1;
		diff_a <= r - b;
		diff_b <= g - b;
	end
	else if (b_ge_r & b_ge_g & r_ge_g) begin
		// B R G
		hue_ofs <= 4'ha;
		diff_a <= r - g;
		diff_b <= b - g;	
	end
	else if (b_ge_r & b_ge_g & g_ge_r) begin
		// B G R
		hue_ofs <= 4'ha;
		sub <= 1'b1;
		diff_a <= g - r;
		diff_b <= b - r;
	end
	else begin
		// R B G
		hue_ofs <= 4'hf;
		sub <= 1'b1;
		diff_a <= b - g;
		diff_b <= r - g;
	end	
end

reg [5:0] hue_tab;

// do some cheap auto scaling to tighten the error bar
reg [11:0] index;
always @(posedge clk) begin
	index <= (diff_a[7] | diff_b[7]) ? {diff_a[7:2],diff_b[7:2]} :
			 (diff_a[6] | diff_b[6]) ? {diff_a[6:1],diff_b[6:1]} :
			 {diff_a[5:0],diff_b[5:0]};
end

always @(posedge clk) begin
	case (index)
			12'd0 : hue_tab <= 6'd0;
			12'd1 : hue_tab <= 6'd0;
			12'd2 : hue_tab <= 6'd0;
			12'd3 : hue_tab <= 6'd0;
			12'd4 : hue_tab <= 6'd0;
			12'd5 : hue_tab <= 6'd0;
			12'd6 : hue_tab <= 6'd0;
			12'd7 : hue_tab <= 6'd0;
			12'd8 : hue_tab <= 6'd0;
			12'd9 : hue_tab <= 6'd0;
			12'd10 : hue_tab <= 6'd0;
			12'd11 : hue_tab <= 6'd0;
			12'd12 : hue_tab <= 6'd0;
			12'd13 : hue_tab <= 6'd0;
			12'd14 : hue_tab <= 6'd0;
			12'd15 : hue_tab <= 6'd0;
			12'd16 : hue_tab <= 6'd0;
			12'd17 : hue_tab <= 6'd0;
			12'd18 : hue_tab <= 6'd0;
			12'd19 : hue_tab <= 6'd0;
			12'd20 : hue_tab <= 6'd0;
			12'd21 : hue_tab <= 6'd0;
			12'd22 : hue_tab <= 6'd0;
			12'd23 : hue_tab <= 6'd0;
			12'd24 : hue_tab <= 6'd0;
			12'd25 : hue_tab <= 6'd0;
			12'd26 : hue_tab <= 6'd0;
			12'd27 : hue_tab <= 6'd0;
			12'd28 : hue_tab <= 6'd0;
			12'd29 : hue_tab <= 6'd0;
			12'd30 : hue_tab <= 6'd0;
			12'd31 : hue_tab <= 6'd0;
			12'd32 : hue_tab <= 6'd0;
			12'd33 : hue_tab <= 6'd0;
			12'd34 : hue_tab <= 6'd0;
			12'd35 : hue_tab <= 6'd0;
			12'd36 : hue_tab <= 6'd0;
			12'd37 : hue_tab <= 6'd0;
			12'd38 : hue_tab <= 6'd0;
			12'd39 : hue_tab <= 6'd0;
			12'd40 : hue_tab <= 6'd0;
			12'd41 : hue_tab <= 6'd0;
			12'd42 : hue_tab <= 6'd0;
			12'd43 : hue_tab <= 6'd0;
			12'd44 : hue_tab <= 6'd0;
			12'd45 : hue_tab <= 6'd0;
			12'd46 : hue_tab <= 6'd0;
			12'd47 : hue_tab <= 6'd0;
			12'd48 : hue_tab <= 6'd0;
			12'd49 : hue_tab <= 6'd0;
			12'd50 : hue_tab <= 6'd0;
			12'd51 : hue_tab <= 6'd0;
			12'd52 : hue_tab <= 6'd0;
			12'd53 : hue_tab <= 6'd0;
			12'd54 : hue_tab <= 6'd0;
			12'd55 : hue_tab <= 6'd0;
			12'd56 : hue_tab <= 6'd0;
			12'd57 : hue_tab <= 6'd0;
			12'd58 : hue_tab <= 6'd0;
			12'd59 : hue_tab <= 6'd0;
			12'd60 : hue_tab <= 6'd0;
			12'd61 : hue_tab <= 6'd0;
			12'd62 : hue_tab <= 6'd0;
			12'd63 : hue_tab <= 6'd0;
			12'd64 : hue_tab <= 6'd0;
			12'd65 : hue_tab <= 6'd40;
			12'd66 : hue_tab <= 6'd20;
			12'd67 : hue_tab <= 6'd13;
			12'd68 : hue_tab <= 6'd10;
			12'd69 : hue_tab <= 6'd8;
			12'd70 : hue_tab <= 6'd6;
			12'd71 : hue_tab <= 6'd5;
			12'd72 : hue_tab <= 6'd5;
			12'd73 : hue_tab <= 6'd4;
			12'd74 : hue_tab <= 6'd4;
			12'd75 : hue_tab <= 6'd3;
			12'd76 : hue_tab <= 6'd3;
			12'd77 : hue_tab <= 6'd3;
			12'd78 : hue_tab <= 6'd2;
			12'd79 : hue_tab <= 6'd2;
			12'd80 : hue_tab <= 6'd2;
			12'd81 : hue_tab <= 6'd2;
			12'd82 : hue_tab <= 6'd2;
			12'd83 : hue_tab <= 6'd2;
			12'd84 : hue_tab <= 6'd2;
			12'd85 : hue_tab <= 6'd1;
			12'd86 : hue_tab <= 6'd1;
			12'd87 : hue_tab <= 6'd1;
			12'd88 : hue_tab <= 6'd1;
			12'd89 : hue_tab <= 6'd1;
			12'd90 : hue_tab <= 6'd1;
			12'd91 : hue_tab <= 6'd1;
			12'd92 : hue_tab <= 6'd1;
			12'd93 : hue_tab <= 6'd1;
			12'd94 : hue_tab <= 6'd1;
			12'd95 : hue_tab <= 6'd1;
			12'd96 : hue_tab <= 6'd1;
			12'd97 : hue_tab <= 6'd1;
			12'd98 : hue_tab <= 6'd1;
			12'd99 : hue_tab <= 6'd1;
			12'd100 : hue_tab <= 6'd1;
			12'd101 : hue_tab <= 6'd1;
			12'd102 : hue_tab <= 6'd1;
			12'd103 : hue_tab <= 6'd1;
			12'd104 : hue_tab <= 6'd1;
			12'd105 : hue_tab <= 6'd0;
			12'd106 : hue_tab <= 6'd0;
			12'd107 : hue_tab <= 6'd0;
			12'd108 : hue_tab <= 6'd0;
			12'd109 : hue_tab <= 6'd0;
			12'd110 : hue_tab <= 6'd0;
			12'd111 : hue_tab <= 6'd0;
			12'd112 : hue_tab <= 6'd0;
			12'd113 : hue_tab <= 6'd0;
			12'd114 : hue_tab <= 6'd0;
			12'd115 : hue_tab <= 6'd0;
			12'd116 : hue_tab <= 6'd0;
			12'd117 : hue_tab <= 6'd0;
			12'd118 : hue_tab <= 6'd0;
			12'd119 : hue_tab <= 6'd0;
			12'd120 : hue_tab <= 6'd0;
			12'd121 : hue_tab <= 6'd0;
			12'd122 : hue_tab <= 6'd0;
			12'd123 : hue_tab <= 6'd0;
			12'd124 : hue_tab <= 6'd0;
			12'd125 : hue_tab <= 6'd0;
			12'd126 : hue_tab <= 6'd0;
			12'd127 : hue_tab <= 6'd0;
			12'd128 : hue_tab <= 6'd0;
			12'd129 : hue_tab <= 6'd40;
			12'd130 : hue_tab <= 6'd40;
			12'd131 : hue_tab <= 6'd26;
			12'd132 : hue_tab <= 6'd20;
			12'd133 : hue_tab <= 6'd16;
			12'd134 : hue_tab <= 6'd13;
			12'd135 : hue_tab <= 6'd11;
			12'd136 : hue_tab <= 6'd10;
			12'd137 : hue_tab <= 6'd8;
			12'd138 : hue_tab <= 6'd8;
			12'd139 : hue_tab <= 6'd7;
			12'd140 : hue_tab <= 6'd6;
			12'd141 : hue_tab <= 6'd6;
			12'd142 : hue_tab <= 6'd5;
			12'd143 : hue_tab <= 6'd5;
			12'd144 : hue_tab <= 6'd5;
			12'd145 : hue_tab <= 6'd4;
			12'd146 : hue_tab <= 6'd4;
			12'd147 : hue_tab <= 6'd4;
			12'd148 : hue_tab <= 6'd4;
			12'd149 : hue_tab <= 6'd3;
			12'd150 : hue_tab <= 6'd3;
			12'd151 : hue_tab <= 6'd3;
			12'd152 : hue_tab <= 6'd3;
			12'd153 : hue_tab <= 6'd3;
			12'd154 : hue_tab <= 6'd3;
			12'd155 : hue_tab <= 6'd2;
			12'd156 : hue_tab <= 6'd2;
			12'd157 : hue_tab <= 6'd2;
			12'd158 : hue_tab <= 6'd2;
			12'd159 : hue_tab <= 6'd2;
			12'd160 : hue_tab <= 6'd2;
			12'd161 : hue_tab <= 6'd2;
			12'd162 : hue_tab <= 6'd2;
			12'd163 : hue_tab <= 6'd2;
			12'd164 : hue_tab <= 6'd2;
			12'd165 : hue_tab <= 6'd2;
			12'd166 : hue_tab <= 6'd2;
			12'd167 : hue_tab <= 6'd2;
			12'd168 : hue_tab <= 6'd2;
			12'd169 : hue_tab <= 6'd1;
			12'd170 : hue_tab <= 6'd1;
			12'd171 : hue_tab <= 6'd1;
			12'd172 : hue_tab <= 6'd1;
			12'd173 : hue_tab <= 6'd1;
			12'd174 : hue_tab <= 6'd1;
			12'd175 : hue_tab <= 6'd1;
			12'd176 : hue_tab <= 6'd1;
			12'd177 : hue_tab <= 6'd1;
			12'd178 : hue_tab <= 6'd1;
			12'd179 : hue_tab <= 6'd1;
			12'd180 : hue_tab <= 6'd1;
			12'd181 : hue_tab <= 6'd1;
			12'd182 : hue_tab <= 6'd1;
			12'd183 : hue_tab <= 6'd1;
			12'd184 : hue_tab <= 6'd1;
			12'd185 : hue_tab <= 6'd1;
			12'd186 : hue_tab <= 6'd1;
			12'd187 : hue_tab <= 6'd1;
			12'd188 : hue_tab <= 6'd1;
			12'd189 : hue_tab <= 6'd1;
			12'd190 : hue_tab <= 6'd1;
			12'd191 : hue_tab <= 6'd1;
			12'd192 : hue_tab <= 6'd0;
			12'd193 : hue_tab <= 6'd40;
			12'd194 : hue_tab <= 6'd40;
			12'd195 : hue_tab <= 6'd40;
			12'd196 : hue_tab <= 6'd30;
			12'd197 : hue_tab <= 6'd24;
			12'd198 : hue_tab <= 6'd20;
			12'd199 : hue_tab <= 6'd17;
			12'd200 : hue_tab <= 6'd15;
			12'd201 : hue_tab <= 6'd13;
			12'd202 : hue_tab <= 6'd12;
			12'd203 : hue_tab <= 6'd10;
			12'd204 : hue_tab <= 6'd10;
			12'd205 : hue_tab <= 6'd9;
			12'd206 : hue_tab <= 6'd8;
			12'd207 : hue_tab <= 6'd8;
			12'd208 : hue_tab <= 6'd7;
			12'd209 : hue_tab <= 6'd7;
			12'd210 : hue_tab <= 6'd6;
			12'd211 : hue_tab <= 6'd6;
			12'd212 : hue_tab <= 6'd6;
			12'd213 : hue_tab <= 6'd5;
			12'd214 : hue_tab <= 6'd5;
			12'd215 : hue_tab <= 6'd5;
			12'd216 : hue_tab <= 6'd5;
			12'd217 : hue_tab <= 6'd4;
			12'd218 : hue_tab <= 6'd4;
			12'd219 : hue_tab <= 6'd4;
			12'd220 : hue_tab <= 6'd4;
			12'd221 : hue_tab <= 6'd4;
			12'd222 : hue_tab <= 6'd4;
			12'd223 : hue_tab <= 6'd3;
			12'd224 : hue_tab <= 6'd3;
			12'd225 : hue_tab <= 6'd3;
			12'd226 : hue_tab <= 6'd3;
			12'd227 : hue_tab <= 6'd3;
			12'd228 : hue_tab <= 6'd3;
			12'd229 : hue_tab <= 6'd3;
			12'd230 : hue_tab <= 6'd3;
			12'd231 : hue_tab <= 6'd3;
			12'd232 : hue_tab <= 6'd3;
			12'd233 : hue_tab <= 6'd2;
			12'd234 : hue_tab <= 6'd2;
			12'd235 : hue_tab <= 6'd2;
			12'd236 : hue_tab <= 6'd2;
			12'd237 : hue_tab <= 6'd2;
			12'd238 : hue_tab <= 6'd2;
			12'd239 : hue_tab <= 6'd2;
			12'd240 : hue_tab <= 6'd2;
			12'd241 : hue_tab <= 6'd2;
			12'd242 : hue_tab <= 6'd2;
			12'd243 : hue_tab <= 6'd2;
			12'd244 : hue_tab <= 6'd2;
			12'd245 : hue_tab <= 6'd2;
			12'd246 : hue_tab <= 6'd2;
			12'd247 : hue_tab <= 6'd2;
			12'd248 : hue_tab <= 6'd2;
			12'd249 : hue_tab <= 6'd2;
			12'd250 : hue_tab <= 6'd2;
			12'd251 : hue_tab <= 6'd2;
			12'd252 : hue_tab <= 6'd2;
			12'd253 : hue_tab <= 6'd1;
			12'd254 : hue_tab <= 6'd1;
			12'd255 : hue_tab <= 6'd1;
			12'd256 : hue_tab <= 6'd0;
			12'd257 : hue_tab <= 6'd40;
			12'd258 : hue_tab <= 6'd40;
			12'd259 : hue_tab <= 6'd40;
			12'd260 : hue_tab <= 6'd40;
			12'd261 : hue_tab <= 6'd32;
			12'd262 : hue_tab <= 6'd26;
			12'd263 : hue_tab <= 6'd22;
			12'd264 : hue_tab <= 6'd20;
			12'd265 : hue_tab <= 6'd17;
			12'd266 : hue_tab <= 6'd16;
			12'd267 : hue_tab <= 6'd14;
			12'd268 : hue_tab <= 6'd13;
			12'd269 : hue_tab <= 6'd12;
			12'd270 : hue_tab <= 6'd11;
			12'd271 : hue_tab <= 6'd10;
			12'd272 : hue_tab <= 6'd10;
			12'd273 : hue_tab <= 6'd9;
			12'd274 : hue_tab <= 6'd8;
			12'd275 : hue_tab <= 6'd8;
			12'd276 : hue_tab <= 6'd8;
			12'd277 : hue_tab <= 6'd7;
			12'd278 : hue_tab <= 6'd7;
			12'd279 : hue_tab <= 6'd6;
			12'd280 : hue_tab <= 6'd6;
			12'd281 : hue_tab <= 6'd6;
			12'd282 : hue_tab <= 6'd6;
			12'd283 : hue_tab <= 6'd5;
			12'd284 : hue_tab <= 6'd5;
			12'd285 : hue_tab <= 6'd5;
			12'd286 : hue_tab <= 6'd5;
			12'd287 : hue_tab <= 6'd5;
			12'd288 : hue_tab <= 6'd5;
			12'd289 : hue_tab <= 6'd4;
			12'd290 : hue_tab <= 6'd4;
			12'd291 : hue_tab <= 6'd4;
			12'd292 : hue_tab <= 6'd4;
			12'd293 : hue_tab <= 6'd4;
			12'd294 : hue_tab <= 6'd4;
			12'd295 : hue_tab <= 6'd4;
			12'd296 : hue_tab <= 6'd4;
			12'd297 : hue_tab <= 6'd3;
			12'd298 : hue_tab <= 6'd3;
			12'd299 : hue_tab <= 6'd3;
			12'd300 : hue_tab <= 6'd3;
			12'd301 : hue_tab <= 6'd3;
			12'd302 : hue_tab <= 6'd3;
			12'd303 : hue_tab <= 6'd3;
			12'd304 : hue_tab <= 6'd3;
			12'd305 : hue_tab <= 6'd3;
			12'd306 : hue_tab <= 6'd3;
			12'd307 : hue_tab <= 6'd3;
			12'd308 : hue_tab <= 6'd3;
			12'd309 : hue_tab <= 6'd3;
			12'd310 : hue_tab <= 6'd2;
			12'd311 : hue_tab <= 6'd2;
			12'd312 : hue_tab <= 6'd2;
			12'd313 : hue_tab <= 6'd2;
			12'd314 : hue_tab <= 6'd2;
			12'd315 : hue_tab <= 6'd2;
			12'd316 : hue_tab <= 6'd2;
			12'd317 : hue_tab <= 6'd2;
			12'd318 : hue_tab <= 6'd2;
			12'd319 : hue_tab <= 6'd2;
			12'd320 : hue_tab <= 6'd0;
			12'd321 : hue_tab <= 6'd40;
			12'd322 : hue_tab <= 6'd40;
			12'd323 : hue_tab <= 6'd40;
			12'd324 : hue_tab <= 6'd40;
			12'd325 : hue_tab <= 6'd40;
			12'd326 : hue_tab <= 6'd33;
			12'd327 : hue_tab <= 6'd28;
			12'd328 : hue_tab <= 6'd25;
			12'd329 : hue_tab <= 6'd22;
			12'd330 : hue_tab <= 6'd20;
			12'd331 : hue_tab <= 6'd18;
			12'd332 : hue_tab <= 6'd16;
			12'd333 : hue_tab <= 6'd15;
			12'd334 : hue_tab <= 6'd14;
			12'd335 : hue_tab <= 6'd13;
			12'd336 : hue_tab <= 6'd12;
			12'd337 : hue_tab <= 6'd11;
			12'd338 : hue_tab <= 6'd11;
			12'd339 : hue_tab <= 6'd10;
			12'd340 : hue_tab <= 6'd10;
			12'd341 : hue_tab <= 6'd9;
			12'd342 : hue_tab <= 6'd9;
			12'd343 : hue_tab <= 6'd8;
			12'd344 : hue_tab <= 6'd8;
			12'd345 : hue_tab <= 6'd8;
			12'd346 : hue_tab <= 6'd7;
			12'd347 : hue_tab <= 6'd7;
			12'd348 : hue_tab <= 6'd7;
			12'd349 : hue_tab <= 6'd6;
			12'd350 : hue_tab <= 6'd6;
			12'd351 : hue_tab <= 6'd6;
			12'd352 : hue_tab <= 6'd6;
			12'd353 : hue_tab <= 6'd6;
			12'd354 : hue_tab <= 6'd5;
			12'd355 : hue_tab <= 6'd5;
			12'd356 : hue_tab <= 6'd5;
			12'd357 : hue_tab <= 6'd5;
			12'd358 : hue_tab <= 6'd5;
			12'd359 : hue_tab <= 6'd5;
			12'd360 : hue_tab <= 6'd5;
			12'd361 : hue_tab <= 6'd4;
			12'd362 : hue_tab <= 6'd4;
			12'd363 : hue_tab <= 6'd4;
			12'd364 : hue_tab <= 6'd4;
			12'd365 : hue_tab <= 6'd4;
			12'd366 : hue_tab <= 6'd4;
			12'd367 : hue_tab <= 6'd4;
			12'd368 : hue_tab <= 6'd4;
			12'd369 : hue_tab <= 6'd4;
			12'd370 : hue_tab <= 6'd4;
			12'd371 : hue_tab <= 6'd3;
			12'd372 : hue_tab <= 6'd3;
			12'd373 : hue_tab <= 6'd3;
			12'd374 : hue_tab <= 6'd3;
			12'd375 : hue_tab <= 6'd3;
			12'd376 : hue_tab <= 6'd3;
			12'd377 : hue_tab <= 6'd3;
			12'd378 : hue_tab <= 6'd3;
			12'd379 : hue_tab <= 6'd3;
			12'd380 : hue_tab <= 6'd3;
			12'd381 : hue_tab <= 6'd3;
			12'd382 : hue_tab <= 6'd3;
			12'd383 : hue_tab <= 6'd3;
			12'd384 : hue_tab <= 6'd0;
			12'd385 : hue_tab <= 6'd40;
			12'd386 : hue_tab <= 6'd40;
			12'd387 : hue_tab <= 6'd40;
			12'd388 : hue_tab <= 6'd40;
			12'd389 : hue_tab <= 6'd40;
			12'd390 : hue_tab <= 6'd40;
			12'd391 : hue_tab <= 6'd34;
			12'd392 : hue_tab <= 6'd30;
			12'd393 : hue_tab <= 6'd26;
			12'd394 : hue_tab <= 6'd24;
			12'd395 : hue_tab <= 6'd21;
			12'd396 : hue_tab <= 6'd20;
			12'd397 : hue_tab <= 6'd18;
			12'd398 : hue_tab <= 6'd17;
			12'd399 : hue_tab <= 6'd16;
			12'd400 : hue_tab <= 6'd15;
			12'd401 : hue_tab <= 6'd14;
			12'd402 : hue_tab <= 6'd13;
			12'd403 : hue_tab <= 6'd12;
			12'd404 : hue_tab <= 6'd12;
			12'd405 : hue_tab <= 6'd11;
			12'd406 : hue_tab <= 6'd10;
			12'd407 : hue_tab <= 6'd10;
			12'd408 : hue_tab <= 6'd10;
			12'd409 : hue_tab <= 6'd9;
			12'd410 : hue_tab <= 6'd9;
			12'd411 : hue_tab <= 6'd8;
			12'd412 : hue_tab <= 6'd8;
			12'd413 : hue_tab <= 6'd8;
			12'd414 : hue_tab <= 6'd8;
			12'd415 : hue_tab <= 6'd7;
			12'd416 : hue_tab <= 6'd7;
			12'd417 : hue_tab <= 6'd7;
			12'd418 : hue_tab <= 6'd7;
			12'd419 : hue_tab <= 6'd6;
			12'd420 : hue_tab <= 6'd6;
			12'd421 : hue_tab <= 6'd6;
			12'd422 : hue_tab <= 6'd6;
			12'd423 : hue_tab <= 6'd6;
			12'd424 : hue_tab <= 6'd6;
			12'd425 : hue_tab <= 6'd5;
			12'd426 : hue_tab <= 6'd5;
			12'd427 : hue_tab <= 6'd5;
			12'd428 : hue_tab <= 6'd5;
			12'd429 : hue_tab <= 6'd5;
			12'd430 : hue_tab <= 6'd5;
			12'd431 : hue_tab <= 6'd5;
			12'd432 : hue_tab <= 6'd5;
			12'd433 : hue_tab <= 6'd4;
			12'd434 : hue_tab <= 6'd4;
			12'd435 : hue_tab <= 6'd4;
			12'd436 : hue_tab <= 6'd4;
			12'd437 : hue_tab <= 6'd4;
			12'd438 : hue_tab <= 6'd4;
			12'd439 : hue_tab <= 6'd4;
			12'd440 : hue_tab <= 6'd4;
			12'd441 : hue_tab <= 6'd4;
			12'd442 : hue_tab <= 6'd4;
			12'd443 : hue_tab <= 6'd4;
			12'd444 : hue_tab <= 6'd4;
			12'd445 : hue_tab <= 6'd3;
			12'd446 : hue_tab <= 6'd3;
			12'd447 : hue_tab <= 6'd3;
			12'd448 : hue_tab <= 6'd0;
			12'd449 : hue_tab <= 6'd40;
			12'd450 : hue_tab <= 6'd40;
			12'd451 : hue_tab <= 6'd40;
			12'd452 : hue_tab <= 6'd40;
			12'd453 : hue_tab <= 6'd40;
			12'd454 : hue_tab <= 6'd40;
			12'd455 : hue_tab <= 6'd40;
			12'd456 : hue_tab <= 6'd35;
			12'd457 : hue_tab <= 6'd31;
			12'd458 : hue_tab <= 6'd28;
			12'd459 : hue_tab <= 6'd25;
			12'd460 : hue_tab <= 6'd23;
			12'd461 : hue_tab <= 6'd21;
			12'd462 : hue_tab <= 6'd20;
			12'd463 : hue_tab <= 6'd18;
			12'd464 : hue_tab <= 6'd17;
			12'd465 : hue_tab <= 6'd16;
			12'd466 : hue_tab <= 6'd15;
			12'd467 : hue_tab <= 6'd14;
			12'd468 : hue_tab <= 6'd14;
			12'd469 : hue_tab <= 6'd13;
			12'd470 : hue_tab <= 6'd12;
			12'd471 : hue_tab <= 6'd12;
			12'd472 : hue_tab <= 6'd11;
			12'd473 : hue_tab <= 6'd11;
			12'd474 : hue_tab <= 6'd10;
			12'd475 : hue_tab <= 6'd10;
			12'd476 : hue_tab <= 6'd10;
			12'd477 : hue_tab <= 6'd9;
			12'd478 : hue_tab <= 6'd9;
			12'd479 : hue_tab <= 6'd9;
			12'd480 : hue_tab <= 6'd8;
			12'd481 : hue_tab <= 6'd8;
			12'd482 : hue_tab <= 6'd8;
			12'd483 : hue_tab <= 6'd8;
			12'd484 : hue_tab <= 6'd7;
			12'd485 : hue_tab <= 6'd7;
			12'd486 : hue_tab <= 6'd7;
			12'd487 : hue_tab <= 6'd7;
			12'd488 : hue_tab <= 6'd7;
			12'd489 : hue_tab <= 6'd6;
			12'd490 : hue_tab <= 6'd6;
			12'd491 : hue_tab <= 6'd6;
			12'd492 : hue_tab <= 6'd6;
			12'd493 : hue_tab <= 6'd6;
			12'd494 : hue_tab <= 6'd6;
			12'd495 : hue_tab <= 6'd5;
			12'd496 : hue_tab <= 6'd5;
			12'd497 : hue_tab <= 6'd5;
			12'd498 : hue_tab <= 6'd5;
			12'd499 : hue_tab <= 6'd5;
			12'd500 : hue_tab <= 6'd5;
			12'd501 : hue_tab <= 6'd5;
			12'd502 : hue_tab <= 6'd5;
			12'd503 : hue_tab <= 6'd5;
			12'd504 : hue_tab <= 6'd5;
			12'd505 : hue_tab <= 6'd4;
			12'd506 : hue_tab <= 6'd4;
			12'd507 : hue_tab <= 6'd4;
			12'd508 : hue_tab <= 6'd4;
			12'd509 : hue_tab <= 6'd4;
			12'd510 : hue_tab <= 6'd4;
			12'd511 : hue_tab <= 6'd4;
			12'd512 : hue_tab <= 6'd0;
			12'd513 : hue_tab <= 6'd40;
			12'd514 : hue_tab <= 6'd40;
			12'd515 : hue_tab <= 6'd40;
			12'd516 : hue_tab <= 6'd40;
			12'd517 : hue_tab <= 6'd40;
			12'd518 : hue_tab <= 6'd40;
			12'd519 : hue_tab <= 6'd40;
			12'd520 : hue_tab <= 6'd40;
			12'd521 : hue_tab <= 6'd35;
			12'd522 : hue_tab <= 6'd32;
			12'd523 : hue_tab <= 6'd29;
			12'd524 : hue_tab <= 6'd26;
			12'd525 : hue_tab <= 6'd24;
			12'd526 : hue_tab <= 6'd22;
			12'd527 : hue_tab <= 6'd21;
			12'd528 : hue_tab <= 6'd20;
			12'd529 : hue_tab <= 6'd18;
			12'd530 : hue_tab <= 6'd17;
			12'd531 : hue_tab <= 6'd16;
			12'd532 : hue_tab <= 6'd16;
			12'd533 : hue_tab <= 6'd15;
			12'd534 : hue_tab <= 6'd14;
			12'd535 : hue_tab <= 6'd13;
			12'd536 : hue_tab <= 6'd13;
			12'd537 : hue_tab <= 6'd12;
			12'd538 : hue_tab <= 6'd12;
			12'd539 : hue_tab <= 6'd11;
			12'd540 : hue_tab <= 6'd11;
			12'd541 : hue_tab <= 6'd11;
			12'd542 : hue_tab <= 6'd10;
			12'd543 : hue_tab <= 6'd10;
			12'd544 : hue_tab <= 6'd10;
			12'd545 : hue_tab <= 6'd9;
			12'd546 : hue_tab <= 6'd9;
			12'd547 : hue_tab <= 6'd9;
			12'd548 : hue_tab <= 6'd8;
			12'd549 : hue_tab <= 6'd8;
			12'd550 : hue_tab <= 6'd8;
			12'd551 : hue_tab <= 6'd8;
			12'd552 : hue_tab <= 6'd8;
			12'd553 : hue_tab <= 6'd7;
			12'd554 : hue_tab <= 6'd7;
			12'd555 : hue_tab <= 6'd7;
			12'd556 : hue_tab <= 6'd7;
			12'd557 : hue_tab <= 6'd7;
			12'd558 : hue_tab <= 6'd6;
			12'd559 : hue_tab <= 6'd6;
			12'd560 : hue_tab <= 6'd6;
			12'd561 : hue_tab <= 6'd6;
			12'd562 : hue_tab <= 6'd6;
			12'd563 : hue_tab <= 6'd6;
			12'd564 : hue_tab <= 6'd6;
			12'd565 : hue_tab <= 6'd6;
			12'd566 : hue_tab <= 6'd5;
			12'd567 : hue_tab <= 6'd5;
			12'd568 : hue_tab <= 6'd5;
			12'd569 : hue_tab <= 6'd5;
			12'd570 : hue_tab <= 6'd5;
			12'd571 : hue_tab <= 6'd5;
			12'd572 : hue_tab <= 6'd5;
			12'd573 : hue_tab <= 6'd5;
			12'd574 : hue_tab <= 6'd5;
			12'd575 : hue_tab <= 6'd5;
			12'd576 : hue_tab <= 6'd0;
			12'd577 : hue_tab <= 6'd40;
			12'd578 : hue_tab <= 6'd40;
			12'd579 : hue_tab <= 6'd40;
			12'd580 : hue_tab <= 6'd40;
			12'd581 : hue_tab <= 6'd40;
			12'd582 : hue_tab <= 6'd40;
			12'd583 : hue_tab <= 6'd40;
			12'd584 : hue_tab <= 6'd40;
			12'd585 : hue_tab <= 6'd40;
			12'd586 : hue_tab <= 6'd36;
			12'd587 : hue_tab <= 6'd32;
			12'd588 : hue_tab <= 6'd30;
			12'd589 : hue_tab <= 6'd27;
			12'd590 : hue_tab <= 6'd25;
			12'd591 : hue_tab <= 6'd24;
			12'd592 : hue_tab <= 6'd22;
			12'd593 : hue_tab <= 6'd21;
			12'd594 : hue_tab <= 6'd20;
			12'd595 : hue_tab <= 6'd18;
			12'd596 : hue_tab <= 6'd18;
			12'd597 : hue_tab <= 6'd17;
			12'd598 : hue_tab <= 6'd16;
			12'd599 : hue_tab <= 6'd15;
			12'd600 : hue_tab <= 6'd15;
			12'd601 : hue_tab <= 6'd14;
			12'd602 : hue_tab <= 6'd13;
			12'd603 : hue_tab <= 6'd13;
			12'd604 : hue_tab <= 6'd12;
			12'd605 : hue_tab <= 6'd12;
			12'd606 : hue_tab <= 6'd12;
			12'd607 : hue_tab <= 6'd11;
			12'd608 : hue_tab <= 6'd11;
			12'd609 : hue_tab <= 6'd10;
			12'd610 : hue_tab <= 6'd10;
			12'd611 : hue_tab <= 6'd10;
			12'd612 : hue_tab <= 6'd10;
			12'd613 : hue_tab <= 6'd9;
			12'd614 : hue_tab <= 6'd9;
			12'd615 : hue_tab <= 6'd9;
			12'd616 : hue_tab <= 6'd9;
			12'd617 : hue_tab <= 6'd8;
			12'd618 : hue_tab <= 6'd8;
			12'd619 : hue_tab <= 6'd8;
			12'd620 : hue_tab <= 6'd8;
			12'd621 : hue_tab <= 6'd8;
			12'd622 : hue_tab <= 6'd7;
			12'd623 : hue_tab <= 6'd7;
			12'd624 : hue_tab <= 6'd7;
			12'd625 : hue_tab <= 6'd7;
			12'd626 : hue_tab <= 6'd7;
			12'd627 : hue_tab <= 6'd7;
			12'd628 : hue_tab <= 6'd6;
			12'd629 : hue_tab <= 6'd6;
			12'd630 : hue_tab <= 6'd6;
			12'd631 : hue_tab <= 6'd6;
			12'd632 : hue_tab <= 6'd6;
			12'd633 : hue_tab <= 6'd6;
			12'd634 : hue_tab <= 6'd6;
			12'd635 : hue_tab <= 6'd6;
			12'd636 : hue_tab <= 6'd6;
			12'd637 : hue_tab <= 6'd5;
			12'd638 : hue_tab <= 6'd5;
			12'd639 : hue_tab <= 6'd5;
			12'd640 : hue_tab <= 6'd0;
			12'd641 : hue_tab <= 6'd40;
			12'd642 : hue_tab <= 6'd40;
			12'd643 : hue_tab <= 6'd40;
			12'd644 : hue_tab <= 6'd40;
			12'd645 : hue_tab <= 6'd40;
			12'd646 : hue_tab <= 6'd40;
			12'd647 : hue_tab <= 6'd40;
			12'd648 : hue_tab <= 6'd40;
			12'd649 : hue_tab <= 6'd40;
			12'd650 : hue_tab <= 6'd40;
			12'd651 : hue_tab <= 6'd36;
			12'd652 : hue_tab <= 6'd33;
			12'd653 : hue_tab <= 6'd30;
			12'd654 : hue_tab <= 6'd28;
			12'd655 : hue_tab <= 6'd26;
			12'd656 : hue_tab <= 6'd25;
			12'd657 : hue_tab <= 6'd23;
			12'd658 : hue_tab <= 6'd22;
			12'd659 : hue_tab <= 6'd21;
			12'd660 : hue_tab <= 6'd20;
			12'd661 : hue_tab <= 6'd19;
			12'd662 : hue_tab <= 6'd18;
			12'd663 : hue_tab <= 6'd17;
			12'd664 : hue_tab <= 6'd16;
			12'd665 : hue_tab <= 6'd16;
			12'd666 : hue_tab <= 6'd15;
			12'd667 : hue_tab <= 6'd14;
			12'd668 : hue_tab <= 6'd14;
			12'd669 : hue_tab <= 6'd13;
			12'd670 : hue_tab <= 6'd13;
			12'd671 : hue_tab <= 6'd12;
			12'd672 : hue_tab <= 6'd12;
			12'd673 : hue_tab <= 6'd12;
			12'd674 : hue_tab <= 6'd11;
			12'd675 : hue_tab <= 6'd11;
			12'd676 : hue_tab <= 6'd11;
			12'd677 : hue_tab <= 6'd10;
			12'd678 : hue_tab <= 6'd10;
			12'd679 : hue_tab <= 6'd10;
			12'd680 : hue_tab <= 6'd10;
			12'd681 : hue_tab <= 6'd9;
			12'd682 : hue_tab <= 6'd9;
			12'd683 : hue_tab <= 6'd9;
			12'd684 : hue_tab <= 6'd9;
			12'd685 : hue_tab <= 6'd8;
			12'd686 : hue_tab <= 6'd8;
			12'd687 : hue_tab <= 6'd8;
			12'd688 : hue_tab <= 6'd8;
			12'd689 : hue_tab <= 6'd8;
			12'd690 : hue_tab <= 6'd8;
			12'd691 : hue_tab <= 6'd7;
			12'd692 : hue_tab <= 6'd7;
			12'd693 : hue_tab <= 6'd7;
			12'd694 : hue_tab <= 6'd7;
			12'd695 : hue_tab <= 6'd7;
			12'd696 : hue_tab <= 6'd7;
			12'd697 : hue_tab <= 6'd7;
			12'd698 : hue_tab <= 6'd6;
			12'd699 : hue_tab <= 6'd6;
			12'd700 : hue_tab <= 6'd6;
			12'd701 : hue_tab <= 6'd6;
			12'd702 : hue_tab <= 6'd6;
			12'd703 : hue_tab <= 6'd6;
			12'd704 : hue_tab <= 6'd0;
			12'd705 : hue_tab <= 6'd40;
			12'd706 : hue_tab <= 6'd40;
			12'd707 : hue_tab <= 6'd40;
			12'd708 : hue_tab <= 6'd40;
			12'd709 : hue_tab <= 6'd40;
			12'd710 : hue_tab <= 6'd40;
			12'd711 : hue_tab <= 6'd40;
			12'd712 : hue_tab <= 6'd40;
			12'd713 : hue_tab <= 6'd40;
			12'd714 : hue_tab <= 6'd40;
			12'd715 : hue_tab <= 6'd40;
			12'd716 : hue_tab <= 6'd36;
			12'd717 : hue_tab <= 6'd33;
			12'd718 : hue_tab <= 6'd31;
			12'd719 : hue_tab <= 6'd29;
			12'd720 : hue_tab <= 6'd27;
			12'd721 : hue_tab <= 6'd25;
			12'd722 : hue_tab <= 6'd24;
			12'd723 : hue_tab <= 6'd23;
			12'd724 : hue_tab <= 6'd22;
			12'd725 : hue_tab <= 6'd20;
			12'd726 : hue_tab <= 6'd20;
			12'd727 : hue_tab <= 6'd19;
			12'd728 : hue_tab <= 6'd18;
			12'd729 : hue_tab <= 6'd17;
			12'd730 : hue_tab <= 6'd16;
			12'd731 : hue_tab <= 6'd16;
			12'd732 : hue_tab <= 6'd15;
			12'd733 : hue_tab <= 6'd15;
			12'd734 : hue_tab <= 6'd14;
			12'd735 : hue_tab <= 6'd14;
			12'd736 : hue_tab <= 6'd13;
			12'd737 : hue_tab <= 6'd13;
			12'd738 : hue_tab <= 6'd12;
			12'd739 : hue_tab <= 6'd12;
			12'd740 : hue_tab <= 6'd12;
			12'd741 : hue_tab <= 6'd11;
			12'd742 : hue_tab <= 6'd11;
			12'd743 : hue_tab <= 6'd11;
			12'd744 : hue_tab <= 6'd11;
			12'd745 : hue_tab <= 6'd10;
			12'd746 : hue_tab <= 6'd10;
			12'd747 : hue_tab <= 6'd10;
			12'd748 : hue_tab <= 6'd10;
			12'd749 : hue_tab <= 6'd9;
			12'd750 : hue_tab <= 6'd9;
			12'd751 : hue_tab <= 6'd9;
			12'd752 : hue_tab <= 6'd9;
			12'd753 : hue_tab <= 6'd8;
			12'd754 : hue_tab <= 6'd8;
			12'd755 : hue_tab <= 6'd8;
			12'd756 : hue_tab <= 6'd8;
			12'd757 : hue_tab <= 6'd8;
			12'd758 : hue_tab <= 6'd8;
			12'd759 : hue_tab <= 6'd8;
			12'd760 : hue_tab <= 6'd7;
			12'd761 : hue_tab <= 6'd7;
			12'd762 : hue_tab <= 6'd7;
			12'd763 : hue_tab <= 6'd7;
			12'd764 : hue_tab <= 6'd7;
			12'd765 : hue_tab <= 6'd7;
			12'd766 : hue_tab <= 6'd7;
			12'd767 : hue_tab <= 6'd6;
			12'd768 : hue_tab <= 6'd0;
			12'd769 : hue_tab <= 6'd40;
			12'd770 : hue_tab <= 6'd40;
			12'd771 : hue_tab <= 6'd40;
			12'd772 : hue_tab <= 6'd40;
			12'd773 : hue_tab <= 6'd40;
			12'd774 : hue_tab <= 6'd40;
			12'd775 : hue_tab <= 6'd40;
			12'd776 : hue_tab <= 6'd40;
			12'd777 : hue_tab <= 6'd40;
			12'd778 : hue_tab <= 6'd40;
			12'd779 : hue_tab <= 6'd40;
			12'd780 : hue_tab <= 6'd40;
			12'd781 : hue_tab <= 6'd36;
			12'd782 : hue_tab <= 6'd34;
			12'd783 : hue_tab <= 6'd32;
			12'd784 : hue_tab <= 6'd30;
			12'd785 : hue_tab <= 6'd28;
			12'd786 : hue_tab <= 6'd26;
			12'd787 : hue_tab <= 6'd25;
			12'd788 : hue_tab <= 6'd24;
			12'd789 : hue_tab <= 6'd22;
			12'd790 : hue_tab <= 6'd21;
			12'd791 : hue_tab <= 6'd20;
			12'd792 : hue_tab <= 6'd20;
			12'd793 : hue_tab <= 6'd19;
			12'd794 : hue_tab <= 6'd18;
			12'd795 : hue_tab <= 6'd17;
			12'd796 : hue_tab <= 6'd17;
			12'd797 : hue_tab <= 6'd16;
			12'd798 : hue_tab <= 6'd16;
			12'd799 : hue_tab <= 6'd15;
			12'd800 : hue_tab <= 6'd15;
			12'd801 : hue_tab <= 6'd14;
			12'd802 : hue_tab <= 6'd14;
			12'd803 : hue_tab <= 6'd13;
			12'd804 : hue_tab <= 6'd13;
			12'd805 : hue_tab <= 6'd12;
			12'd806 : hue_tab <= 6'd12;
			12'd807 : hue_tab <= 6'd12;
			12'd808 : hue_tab <= 6'd12;
			12'd809 : hue_tab <= 6'd11;
			12'd810 : hue_tab <= 6'd11;
			12'd811 : hue_tab <= 6'd11;
			12'd812 : hue_tab <= 6'd10;
			12'd813 : hue_tab <= 6'd10;
			12'd814 : hue_tab <= 6'd10;
			12'd815 : hue_tab <= 6'd10;
			12'd816 : hue_tab <= 6'd10;
			12'd817 : hue_tab <= 6'd9;
			12'd818 : hue_tab <= 6'd9;
			12'd819 : hue_tab <= 6'd9;
			12'd820 : hue_tab <= 6'd9;
			12'd821 : hue_tab <= 6'd9;
			12'd822 : hue_tab <= 6'd8;
			12'd823 : hue_tab <= 6'd8;
			12'd824 : hue_tab <= 6'd8;
			12'd825 : hue_tab <= 6'd8;
			12'd826 : hue_tab <= 6'd8;
			12'd827 : hue_tab <= 6'd8;
			12'd828 : hue_tab <= 6'd8;
			12'd829 : hue_tab <= 6'd7;
			12'd830 : hue_tab <= 6'd7;
			12'd831 : hue_tab <= 6'd7;
			12'd832 : hue_tab <= 6'd0;
			12'd833 : hue_tab <= 6'd40;
			12'd834 : hue_tab <= 6'd40;
			12'd835 : hue_tab <= 6'd40;
			12'd836 : hue_tab <= 6'd40;
			12'd837 : hue_tab <= 6'd40;
			12'd838 : hue_tab <= 6'd40;
			12'd839 : hue_tab <= 6'd40;
			12'd840 : hue_tab <= 6'd40;
			12'd841 : hue_tab <= 6'd40;
			12'd842 : hue_tab <= 6'd40;
			12'd843 : hue_tab <= 6'd40;
			12'd844 : hue_tab <= 6'd40;
			12'd845 : hue_tab <= 6'd40;
			12'd846 : hue_tab <= 6'd37;
			12'd847 : hue_tab <= 6'd34;
			12'd848 : hue_tab <= 6'd32;
			12'd849 : hue_tab <= 6'd30;
			12'd850 : hue_tab <= 6'd28;
			12'd851 : hue_tab <= 6'd27;
			12'd852 : hue_tab <= 6'd26;
			12'd853 : hue_tab <= 6'd24;
			12'd854 : hue_tab <= 6'd23;
			12'd855 : hue_tab <= 6'd22;
			12'd856 : hue_tab <= 6'd21;
			12'd857 : hue_tab <= 6'd20;
			12'd858 : hue_tab <= 6'd20;
			12'd859 : hue_tab <= 6'd19;
			12'd860 : hue_tab <= 6'd18;
			12'd861 : hue_tab <= 6'd17;
			12'd862 : hue_tab <= 6'd17;
			12'd863 : hue_tab <= 6'd16;
			12'd864 : hue_tab <= 6'd16;
			12'd865 : hue_tab <= 6'd15;
			12'd866 : hue_tab <= 6'd15;
			12'd867 : hue_tab <= 6'd14;
			12'd868 : hue_tab <= 6'd14;
			12'd869 : hue_tab <= 6'd14;
			12'd870 : hue_tab <= 6'd13;
			12'd871 : hue_tab <= 6'd13;
			12'd872 : hue_tab <= 6'd13;
			12'd873 : hue_tab <= 6'd12;
			12'd874 : hue_tab <= 6'd12;
			12'd875 : hue_tab <= 6'd12;
			12'd876 : hue_tab <= 6'd11;
			12'd877 : hue_tab <= 6'd11;
			12'd878 : hue_tab <= 6'd11;
			12'd879 : hue_tab <= 6'd11;
			12'd880 : hue_tab <= 6'd10;
			12'd881 : hue_tab <= 6'd10;
			12'd882 : hue_tab <= 6'd10;
			12'd883 : hue_tab <= 6'd10;
			12'd884 : hue_tab <= 6'd10;
			12'd885 : hue_tab <= 6'd9;
			12'd886 : hue_tab <= 6'd9;
			12'd887 : hue_tab <= 6'd9;
			12'd888 : hue_tab <= 6'd9;
			12'd889 : hue_tab <= 6'd9;
			12'd890 : hue_tab <= 6'd8;
			12'd891 : hue_tab <= 6'd8;
			12'd892 : hue_tab <= 6'd8;
			12'd893 : hue_tab <= 6'd8;
			12'd894 : hue_tab <= 6'd8;
			12'd895 : hue_tab <= 6'd8;
			12'd896 : hue_tab <= 6'd0;
			12'd897 : hue_tab <= 6'd40;
			12'd898 : hue_tab <= 6'd40;
			12'd899 : hue_tab <= 6'd40;
			12'd900 : hue_tab <= 6'd40;
			12'd901 : hue_tab <= 6'd40;
			12'd902 : hue_tab <= 6'd40;
			12'd903 : hue_tab <= 6'd40;
			12'd904 : hue_tab <= 6'd40;
			12'd905 : hue_tab <= 6'd40;
			12'd906 : hue_tab <= 6'd40;
			12'd907 : hue_tab <= 6'd40;
			12'd908 : hue_tab <= 6'd40;
			12'd909 : hue_tab <= 6'd40;
			12'd910 : hue_tab <= 6'd40;
			12'd911 : hue_tab <= 6'd37;
			12'd912 : hue_tab <= 6'd35;
			12'd913 : hue_tab <= 6'd32;
			12'd914 : hue_tab <= 6'd31;
			12'd915 : hue_tab <= 6'd29;
			12'd916 : hue_tab <= 6'd28;
			12'd917 : hue_tab <= 6'd26;
			12'd918 : hue_tab <= 6'd25;
			12'd919 : hue_tab <= 6'd24;
			12'd920 : hue_tab <= 6'd23;
			12'd921 : hue_tab <= 6'd22;
			12'd922 : hue_tab <= 6'd21;
			12'd923 : hue_tab <= 6'd20;
			12'd924 : hue_tab <= 6'd20;
			12'd925 : hue_tab <= 6'd19;
			12'd926 : hue_tab <= 6'd18;
			12'd927 : hue_tab <= 6'd18;
			12'd928 : hue_tab <= 6'd17;
			12'd929 : hue_tab <= 6'd16;
			12'd930 : hue_tab <= 6'd16;
			12'd931 : hue_tab <= 6'd16;
			12'd932 : hue_tab <= 6'd15;
			12'd933 : hue_tab <= 6'd15;
			12'd934 : hue_tab <= 6'd14;
			12'd935 : hue_tab <= 6'd14;
			12'd936 : hue_tab <= 6'd14;
			12'd937 : hue_tab <= 6'd13;
			12'd938 : hue_tab <= 6'd13;
			12'd939 : hue_tab <= 6'd13;
			12'd940 : hue_tab <= 6'd12;
			12'd941 : hue_tab <= 6'd12;
			12'd942 : hue_tab <= 6'd12;
			12'd943 : hue_tab <= 6'd11;
			12'd944 : hue_tab <= 6'd11;
			12'd945 : hue_tab <= 6'd11;
			12'd946 : hue_tab <= 6'd11;
			12'd947 : hue_tab <= 6'd10;
			12'd948 : hue_tab <= 6'd10;
			12'd949 : hue_tab <= 6'd10;
			12'd950 : hue_tab <= 6'd10;
			12'd951 : hue_tab <= 6'd10;
			12'd952 : hue_tab <= 6'd10;
			12'd953 : hue_tab <= 6'd9;
			12'd954 : hue_tab <= 6'd9;
			12'd955 : hue_tab <= 6'd9;
			12'd956 : hue_tab <= 6'd9;
			12'd957 : hue_tab <= 6'd9;
			12'd958 : hue_tab <= 6'd9;
			12'd959 : hue_tab <= 6'd8;
			12'd960 : hue_tab <= 6'd0;
			12'd961 : hue_tab <= 6'd40;
			12'd962 : hue_tab <= 6'd40;
			12'd963 : hue_tab <= 6'd40;
			12'd964 : hue_tab <= 6'd40;
			12'd965 : hue_tab <= 6'd40;
			12'd966 : hue_tab <= 6'd40;
			12'd967 : hue_tab <= 6'd40;
			12'd968 : hue_tab <= 6'd40;
			12'd969 : hue_tab <= 6'd40;
			12'd970 : hue_tab <= 6'd40;
			12'd971 : hue_tab <= 6'd40;
			12'd972 : hue_tab <= 6'd40;
			12'd973 : hue_tab <= 6'd40;
			12'd974 : hue_tab <= 6'd40;
			12'd975 : hue_tab <= 6'd40;
			12'd976 : hue_tab <= 6'd37;
			12'd977 : hue_tab <= 6'd35;
			12'd978 : hue_tab <= 6'd33;
			12'd979 : hue_tab <= 6'd31;
			12'd980 : hue_tab <= 6'd30;
			12'd981 : hue_tab <= 6'd28;
			12'd982 : hue_tab <= 6'd27;
			12'd983 : hue_tab <= 6'd26;
			12'd984 : hue_tab <= 6'd25;
			12'd985 : hue_tab <= 6'd24;
			12'd986 : hue_tab <= 6'd23;
			12'd987 : hue_tab <= 6'd22;
			12'd988 : hue_tab <= 6'd21;
			12'd989 : hue_tab <= 6'd20;
			12'd990 : hue_tab <= 6'd20;
			12'd991 : hue_tab <= 6'd19;
			12'd992 : hue_tab <= 6'd18;
			12'd993 : hue_tab <= 6'd18;
			12'd994 : hue_tab <= 6'd17;
			12'd995 : hue_tab <= 6'd17;
			12'd996 : hue_tab <= 6'd16;
			12'd997 : hue_tab <= 6'd16;
			12'd998 : hue_tab <= 6'd15;
			12'd999 : hue_tab <= 6'd15;
			12'd1000 : hue_tab <= 6'd15;
			12'd1001 : hue_tab <= 6'd14;
			12'd1002 : hue_tab <= 6'd14;
			12'd1003 : hue_tab <= 6'd13;
			12'd1004 : hue_tab <= 6'd13;
			12'd1005 : hue_tab <= 6'd13;
			12'd1006 : hue_tab <= 6'd13;
			12'd1007 : hue_tab <= 6'd12;
			12'd1008 : hue_tab <= 6'd12;
			12'd1009 : hue_tab <= 6'd12;
			12'd1010 : hue_tab <= 6'd12;
			12'd1011 : hue_tab <= 6'd11;
			12'd1012 : hue_tab <= 6'd11;
			12'd1013 : hue_tab <= 6'd11;
			12'd1014 : hue_tab <= 6'd11;
			12'd1015 : hue_tab <= 6'd10;
			12'd1016 : hue_tab <= 6'd10;
			12'd1017 : hue_tab <= 6'd10;
			12'd1018 : hue_tab <= 6'd10;
			12'd1019 : hue_tab <= 6'd10;
			12'd1020 : hue_tab <= 6'd10;
			12'd1021 : hue_tab <= 6'd9;
			12'd1022 : hue_tab <= 6'd9;
			12'd1023 : hue_tab <= 6'd9;
			12'd1024 : hue_tab <= 6'd0;
			12'd1025 : hue_tab <= 6'd40;
			12'd1026 : hue_tab <= 6'd40;
			12'd1027 : hue_tab <= 6'd40;
			12'd1028 : hue_tab <= 6'd40;
			12'd1029 : hue_tab <= 6'd40;
			12'd1030 : hue_tab <= 6'd40;
			12'd1031 : hue_tab <= 6'd40;
			12'd1032 : hue_tab <= 6'd40;
			12'd1033 : hue_tab <= 6'd40;
			12'd1034 : hue_tab <= 6'd40;
			12'd1035 : hue_tab <= 6'd40;
			12'd1036 : hue_tab <= 6'd40;
			12'd1037 : hue_tab <= 6'd40;
			12'd1038 : hue_tab <= 6'd40;
			12'd1039 : hue_tab <= 6'd40;
			12'd1040 : hue_tab <= 6'd40;
			12'd1041 : hue_tab <= 6'd37;
			12'd1042 : hue_tab <= 6'd35;
			12'd1043 : hue_tab <= 6'd33;
			12'd1044 : hue_tab <= 6'd32;
			12'd1045 : hue_tab <= 6'd30;
			12'd1046 : hue_tab <= 6'd29;
			12'd1047 : hue_tab <= 6'd27;
			12'd1048 : hue_tab <= 6'd26;
			12'd1049 : hue_tab <= 6'd25;
			12'd1050 : hue_tab <= 6'd24;
			12'd1051 : hue_tab <= 6'd23;
			12'd1052 : hue_tab <= 6'd22;
			12'd1053 : hue_tab <= 6'd22;
			12'd1054 : hue_tab <= 6'd21;
			12'd1055 : hue_tab <= 6'd20;
			12'd1056 : hue_tab <= 6'd20;
			12'd1057 : hue_tab <= 6'd19;
			12'd1058 : hue_tab <= 6'd18;
			12'd1059 : hue_tab <= 6'd18;
			12'd1060 : hue_tab <= 6'd17;
			12'd1061 : hue_tab <= 6'd17;
			12'd1062 : hue_tab <= 6'd16;
			12'd1063 : hue_tab <= 6'd16;
			12'd1064 : hue_tab <= 6'd16;
			12'd1065 : hue_tab <= 6'd15;
			12'd1066 : hue_tab <= 6'd15;
			12'd1067 : hue_tab <= 6'd14;
			12'd1068 : hue_tab <= 6'd14;
			12'd1069 : hue_tab <= 6'd14;
			12'd1070 : hue_tab <= 6'd13;
			12'd1071 : hue_tab <= 6'd13;
			12'd1072 : hue_tab <= 6'd13;
			12'd1073 : hue_tab <= 6'd13;
			12'd1074 : hue_tab <= 6'd12;
			12'd1075 : hue_tab <= 6'd12;
			12'd1076 : hue_tab <= 6'd12;
			12'd1077 : hue_tab <= 6'd12;
			12'd1078 : hue_tab <= 6'd11;
			12'd1079 : hue_tab <= 6'd11;
			12'd1080 : hue_tab <= 6'd11;
			12'd1081 : hue_tab <= 6'd11;
			12'd1082 : hue_tab <= 6'd11;
			12'd1083 : hue_tab <= 6'd10;
			12'd1084 : hue_tab <= 6'd10;
			12'd1085 : hue_tab <= 6'd10;
			12'd1086 : hue_tab <= 6'd10;
			12'd1087 : hue_tab <= 6'd10;
			12'd1088 : hue_tab <= 6'd0;
			12'd1089 : hue_tab <= 6'd40;
			12'd1090 : hue_tab <= 6'd40;
			12'd1091 : hue_tab <= 6'd40;
			12'd1092 : hue_tab <= 6'd40;
			12'd1093 : hue_tab <= 6'd40;
			12'd1094 : hue_tab <= 6'd40;
			12'd1095 : hue_tab <= 6'd40;
			12'd1096 : hue_tab <= 6'd40;
			12'd1097 : hue_tab <= 6'd40;
			12'd1098 : hue_tab <= 6'd40;
			12'd1099 : hue_tab <= 6'd40;
			12'd1100 : hue_tab <= 6'd40;
			12'd1101 : hue_tab <= 6'd40;
			12'd1102 : hue_tab <= 6'd40;
			12'd1103 : hue_tab <= 6'd40;
			12'd1104 : hue_tab <= 6'd40;
			12'd1105 : hue_tab <= 6'd40;
			12'd1106 : hue_tab <= 6'd37;
			12'd1107 : hue_tab <= 6'd35;
			12'd1108 : hue_tab <= 6'd34;
			12'd1109 : hue_tab <= 6'd32;
			12'd1110 : hue_tab <= 6'd30;
			12'd1111 : hue_tab <= 6'd29;
			12'd1112 : hue_tab <= 6'd28;
			12'd1113 : hue_tab <= 6'd27;
			12'd1114 : hue_tab <= 6'd26;
			12'd1115 : hue_tab <= 6'd25;
			12'd1116 : hue_tab <= 6'd24;
			12'd1117 : hue_tab <= 6'd23;
			12'd1118 : hue_tab <= 6'd22;
			12'd1119 : hue_tab <= 6'd21;
			12'd1120 : hue_tab <= 6'd21;
			12'd1121 : hue_tab <= 6'd20;
			12'd1122 : hue_tab <= 6'd20;
			12'd1123 : hue_tab <= 6'd19;
			12'd1124 : hue_tab <= 6'd18;
			12'd1125 : hue_tab <= 6'd18;
			12'd1126 : hue_tab <= 6'd17;
			12'd1127 : hue_tab <= 6'd17;
			12'd1128 : hue_tab <= 6'd17;
			12'd1129 : hue_tab <= 6'd16;
			12'd1130 : hue_tab <= 6'd16;
			12'd1131 : hue_tab <= 6'd15;
			12'd1132 : hue_tab <= 6'd15;
			12'd1133 : hue_tab <= 6'd15;
			12'd1134 : hue_tab <= 6'd14;
			12'd1135 : hue_tab <= 6'd14;
			12'd1136 : hue_tab <= 6'd14;
			12'd1137 : hue_tab <= 6'd13;
			12'd1138 : hue_tab <= 6'd13;
			12'd1139 : hue_tab <= 6'd13;
			12'd1140 : hue_tab <= 6'd13;
			12'd1141 : hue_tab <= 6'd12;
			12'd1142 : hue_tab <= 6'd12;
			12'd1143 : hue_tab <= 6'd12;
			12'd1144 : hue_tab <= 6'd12;
			12'd1145 : hue_tab <= 6'd11;
			12'd1146 : hue_tab <= 6'd11;
			12'd1147 : hue_tab <= 6'd11;
			12'd1148 : hue_tab <= 6'd11;
			12'd1149 : hue_tab <= 6'd11;
			12'd1150 : hue_tab <= 6'd10;
			12'd1151 : hue_tab <= 6'd10;
			12'd1152 : hue_tab <= 6'd0;
			12'd1153 : hue_tab <= 6'd40;
			12'd1154 : hue_tab <= 6'd40;
			12'd1155 : hue_tab <= 6'd40;
			12'd1156 : hue_tab <= 6'd40;
			12'd1157 : hue_tab <= 6'd40;
			12'd1158 : hue_tab <= 6'd40;
			12'd1159 : hue_tab <= 6'd40;
			12'd1160 : hue_tab <= 6'd40;
			12'd1161 : hue_tab <= 6'd40;
			12'd1162 : hue_tab <= 6'd40;
			12'd1163 : hue_tab <= 6'd40;
			12'd1164 : hue_tab <= 6'd40;
			12'd1165 : hue_tab <= 6'd40;
			12'd1166 : hue_tab <= 6'd40;
			12'd1167 : hue_tab <= 6'd40;
			12'd1168 : hue_tab <= 6'd40;
			12'd1169 : hue_tab <= 6'd40;
			12'd1170 : hue_tab <= 6'd40;
			12'd1171 : hue_tab <= 6'd37;
			12'd1172 : hue_tab <= 6'd36;
			12'd1173 : hue_tab <= 6'd34;
			12'd1174 : hue_tab <= 6'd32;
			12'd1175 : hue_tab <= 6'd31;
			12'd1176 : hue_tab <= 6'd30;
			12'd1177 : hue_tab <= 6'd28;
			12'd1178 : hue_tab <= 6'd27;
			12'd1179 : hue_tab <= 6'd26;
			12'd1180 : hue_tab <= 6'd25;
			12'd1181 : hue_tab <= 6'd24;
			12'd1182 : hue_tab <= 6'd24;
			12'd1183 : hue_tab <= 6'd23;
			12'd1184 : hue_tab <= 6'd22;
			12'd1185 : hue_tab <= 6'd21;
			12'd1186 : hue_tab <= 6'd21;
			12'd1187 : hue_tab <= 6'd20;
			12'd1188 : hue_tab <= 6'd20;
			12'd1189 : hue_tab <= 6'd19;
			12'd1190 : hue_tab <= 6'd18;
			12'd1191 : hue_tab <= 6'd18;
			12'd1192 : hue_tab <= 6'd18;
			12'd1193 : hue_tab <= 6'd17;
			12'd1194 : hue_tab <= 6'd17;
			12'd1195 : hue_tab <= 6'd16;
			12'd1196 : hue_tab <= 6'd16;
			12'd1197 : hue_tab <= 6'd16;
			12'd1198 : hue_tab <= 6'd15;
			12'd1199 : hue_tab <= 6'd15;
			12'd1200 : hue_tab <= 6'd15;
			12'd1201 : hue_tab <= 6'd14;
			12'd1202 : hue_tab <= 6'd14;
			12'd1203 : hue_tab <= 6'd14;
			12'd1204 : hue_tab <= 6'd13;
			12'd1205 : hue_tab <= 6'd13;
			12'd1206 : hue_tab <= 6'd13;
			12'd1207 : hue_tab <= 6'd13;
			12'd1208 : hue_tab <= 6'd12;
			12'd1209 : hue_tab <= 6'd12;
			12'd1210 : hue_tab <= 6'd12;
			12'd1211 : hue_tab <= 6'd12;
			12'd1212 : hue_tab <= 6'd12;
			12'd1213 : hue_tab <= 6'd11;
			12'd1214 : hue_tab <= 6'd11;
			12'd1215 : hue_tab <= 6'd11;
			12'd1216 : hue_tab <= 6'd0;
			12'd1217 : hue_tab <= 6'd40;
			12'd1218 : hue_tab <= 6'd40;
			12'd1219 : hue_tab <= 6'd40;
			12'd1220 : hue_tab <= 6'd40;
			12'd1221 : hue_tab <= 6'd40;
			12'd1222 : hue_tab <= 6'd40;
			12'd1223 : hue_tab <= 6'd40;
			12'd1224 : hue_tab <= 6'd40;
			12'd1225 : hue_tab <= 6'd40;
			12'd1226 : hue_tab <= 6'd40;
			12'd1227 : hue_tab <= 6'd40;
			12'd1228 : hue_tab <= 6'd40;
			12'd1229 : hue_tab <= 6'd40;
			12'd1230 : hue_tab <= 6'd40;
			12'd1231 : hue_tab <= 6'd40;
			12'd1232 : hue_tab <= 6'd40;
			12'd1233 : hue_tab <= 6'd40;
			12'd1234 : hue_tab <= 6'd40;
			12'd1235 : hue_tab <= 6'd40;
			12'd1236 : hue_tab <= 6'd38;
			12'd1237 : hue_tab <= 6'd36;
			12'd1238 : hue_tab <= 6'd34;
			12'd1239 : hue_tab <= 6'd33;
			12'd1240 : hue_tab <= 6'd31;
			12'd1241 : hue_tab <= 6'd30;
			12'd1242 : hue_tab <= 6'd29;
			12'd1243 : hue_tab <= 6'd28;
			12'd1244 : hue_tab <= 6'd27;
			12'd1245 : hue_tab <= 6'd26;
			12'd1246 : hue_tab <= 6'd25;
			12'd1247 : hue_tab <= 6'd24;
			12'd1248 : hue_tab <= 6'd23;
			12'd1249 : hue_tab <= 6'd23;
			12'd1250 : hue_tab <= 6'd22;
			12'd1251 : hue_tab <= 6'd21;
			12'd1252 : hue_tab <= 6'd21;
			12'd1253 : hue_tab <= 6'd20;
			12'd1254 : hue_tab <= 6'd20;
			12'd1255 : hue_tab <= 6'd19;
			12'd1256 : hue_tab <= 6'd19;
			12'd1257 : hue_tab <= 6'd18;
			12'd1258 : hue_tab <= 6'd18;
			12'd1259 : hue_tab <= 6'd17;
			12'd1260 : hue_tab <= 6'd17;
			12'd1261 : hue_tab <= 6'd16;
			12'd1262 : hue_tab <= 6'd16;
			12'd1263 : hue_tab <= 6'd16;
			12'd1264 : hue_tab <= 6'd15;
			12'd1265 : hue_tab <= 6'd15;
			12'd1266 : hue_tab <= 6'd15;
			12'd1267 : hue_tab <= 6'd14;
			12'd1268 : hue_tab <= 6'd14;
			12'd1269 : hue_tab <= 6'd14;
			12'd1270 : hue_tab <= 6'd14;
			12'd1271 : hue_tab <= 6'd13;
			12'd1272 : hue_tab <= 6'd13;
			12'd1273 : hue_tab <= 6'd13;
			12'd1274 : hue_tab <= 6'd13;
			12'd1275 : hue_tab <= 6'd12;
			12'd1276 : hue_tab <= 6'd12;
			12'd1277 : hue_tab <= 6'd12;
			12'd1278 : hue_tab <= 6'd12;
			12'd1279 : hue_tab <= 6'd12;
			12'd1280 : hue_tab <= 6'd0;
			12'd1281 : hue_tab <= 6'd40;
			12'd1282 : hue_tab <= 6'd40;
			12'd1283 : hue_tab <= 6'd40;
			12'd1284 : hue_tab <= 6'd40;
			12'd1285 : hue_tab <= 6'd40;
			12'd1286 : hue_tab <= 6'd40;
			12'd1287 : hue_tab <= 6'd40;
			12'd1288 : hue_tab <= 6'd40;
			12'd1289 : hue_tab <= 6'd40;
			12'd1290 : hue_tab <= 6'd40;
			12'd1291 : hue_tab <= 6'd40;
			12'd1292 : hue_tab <= 6'd40;
			12'd1293 : hue_tab <= 6'd40;
			12'd1294 : hue_tab <= 6'd40;
			12'd1295 : hue_tab <= 6'd40;
			12'd1296 : hue_tab <= 6'd40;
			12'd1297 : hue_tab <= 6'd40;
			12'd1298 : hue_tab <= 6'd40;
			12'd1299 : hue_tab <= 6'd40;
			12'd1300 : hue_tab <= 6'd40;
			12'd1301 : hue_tab <= 6'd38;
			12'd1302 : hue_tab <= 6'd36;
			12'd1303 : hue_tab <= 6'd34;
			12'd1304 : hue_tab <= 6'd33;
			12'd1305 : hue_tab <= 6'd32;
			12'd1306 : hue_tab <= 6'd30;
			12'd1307 : hue_tab <= 6'd29;
			12'd1308 : hue_tab <= 6'd28;
			12'd1309 : hue_tab <= 6'd27;
			12'd1310 : hue_tab <= 6'd26;
			12'd1311 : hue_tab <= 6'd25;
			12'd1312 : hue_tab <= 6'd25;
			12'd1313 : hue_tab <= 6'd24;
			12'd1314 : hue_tab <= 6'd23;
			12'd1315 : hue_tab <= 6'd22;
			12'd1316 : hue_tab <= 6'd22;
			12'd1317 : hue_tab <= 6'd21;
			12'd1318 : hue_tab <= 6'd21;
			12'd1319 : hue_tab <= 6'd20;
			12'd1320 : hue_tab <= 6'd20;
			12'd1321 : hue_tab <= 6'd19;
			12'd1322 : hue_tab <= 6'd19;
			12'd1323 : hue_tab <= 6'd18;
			12'd1324 : hue_tab <= 6'd18;
			12'd1325 : hue_tab <= 6'd17;
			12'd1326 : hue_tab <= 6'd17;
			12'd1327 : hue_tab <= 6'd17;
			12'd1328 : hue_tab <= 6'd16;
			12'd1329 : hue_tab <= 6'd16;
			12'd1330 : hue_tab <= 6'd16;
			12'd1331 : hue_tab <= 6'd15;
			12'd1332 : hue_tab <= 6'd15;
			12'd1333 : hue_tab <= 6'd15;
			12'd1334 : hue_tab <= 6'd14;
			12'd1335 : hue_tab <= 6'd14;
			12'd1336 : hue_tab <= 6'd14;
			12'd1337 : hue_tab <= 6'd14;
			12'd1338 : hue_tab <= 6'd13;
			12'd1339 : hue_tab <= 6'd13;
			12'd1340 : hue_tab <= 6'd13;
			12'd1341 : hue_tab <= 6'd13;
			12'd1342 : hue_tab <= 6'd12;
			12'd1343 : hue_tab <= 6'd12;
			12'd1344 : hue_tab <= 6'd0;
			12'd1345 : hue_tab <= 6'd40;
			12'd1346 : hue_tab <= 6'd40;
			12'd1347 : hue_tab <= 6'd40;
			12'd1348 : hue_tab <= 6'd40;
			12'd1349 : hue_tab <= 6'd40;
			12'd1350 : hue_tab <= 6'd40;
			12'd1351 : hue_tab <= 6'd40;
			12'd1352 : hue_tab <= 6'd40;
			12'd1353 : hue_tab <= 6'd40;
			12'd1354 : hue_tab <= 6'd40;
			12'd1355 : hue_tab <= 6'd40;
			12'd1356 : hue_tab <= 6'd40;
			12'd1357 : hue_tab <= 6'd40;
			12'd1358 : hue_tab <= 6'd40;
			12'd1359 : hue_tab <= 6'd40;
			12'd1360 : hue_tab <= 6'd40;
			12'd1361 : hue_tab <= 6'd40;
			12'd1362 : hue_tab <= 6'd40;
			12'd1363 : hue_tab <= 6'd40;
			12'd1364 : hue_tab <= 6'd40;
			12'd1365 : hue_tab <= 6'd40;
			12'd1366 : hue_tab <= 6'd38;
			12'd1367 : hue_tab <= 6'd36;
			12'd1368 : hue_tab <= 6'd35;
			12'd1369 : hue_tab <= 6'd33;
			12'd1370 : hue_tab <= 6'd32;
			12'd1371 : hue_tab <= 6'd31;
			12'd1372 : hue_tab <= 6'd30;
			12'd1373 : hue_tab <= 6'd28;
			12'd1374 : hue_tab <= 6'd28;
			12'd1375 : hue_tab <= 6'd27;
			12'd1376 : hue_tab <= 6'd26;
			12'd1377 : hue_tab <= 6'd25;
			12'd1378 : hue_tab <= 6'd24;
			12'd1379 : hue_tab <= 6'd24;
			12'd1380 : hue_tab <= 6'd23;
			12'd1381 : hue_tab <= 6'd22;
			12'd1382 : hue_tab <= 6'd22;
			12'd1383 : hue_tab <= 6'd21;
			12'd1384 : hue_tab <= 6'd21;
			12'd1385 : hue_tab <= 6'd20;
			12'd1386 : hue_tab <= 6'd20;
			12'd1387 : hue_tab <= 6'd19;
			12'd1388 : hue_tab <= 6'd19;
			12'd1389 : hue_tab <= 6'd18;
			12'd1390 : hue_tab <= 6'd18;
			12'd1391 : hue_tab <= 6'd17;
			12'd1392 : hue_tab <= 6'd17;
			12'd1393 : hue_tab <= 6'd17;
			12'd1394 : hue_tab <= 6'd16;
			12'd1395 : hue_tab <= 6'd16;
			12'd1396 : hue_tab <= 6'd16;
			12'd1397 : hue_tab <= 6'd15;
			12'd1398 : hue_tab <= 6'd15;
			12'd1399 : hue_tab <= 6'd15;
			12'd1400 : hue_tab <= 6'd15;
			12'd1401 : hue_tab <= 6'd14;
			12'd1402 : hue_tab <= 6'd14;
			12'd1403 : hue_tab <= 6'd14;
			12'd1404 : hue_tab <= 6'd14;
			12'd1405 : hue_tab <= 6'd13;
			12'd1406 : hue_tab <= 6'd13;
			12'd1407 : hue_tab <= 6'd13;
			12'd1408 : hue_tab <= 6'd0;
			12'd1409 : hue_tab <= 6'd40;
			12'd1410 : hue_tab <= 6'd40;
			12'd1411 : hue_tab <= 6'd40;
			12'd1412 : hue_tab <= 6'd40;
			12'd1413 : hue_tab <= 6'd40;
			12'd1414 : hue_tab <= 6'd40;
			12'd1415 : hue_tab <= 6'd40;
			12'd1416 : hue_tab <= 6'd40;
			12'd1417 : hue_tab <= 6'd40;
			12'd1418 : hue_tab <= 6'd40;
			12'd1419 : hue_tab <= 6'd40;
			12'd1420 : hue_tab <= 6'd40;
			12'd1421 : hue_tab <= 6'd40;
			12'd1422 : hue_tab <= 6'd40;
			12'd1423 : hue_tab <= 6'd40;
			12'd1424 : hue_tab <= 6'd40;
			12'd1425 : hue_tab <= 6'd40;
			12'd1426 : hue_tab <= 6'd40;
			12'd1427 : hue_tab <= 6'd40;
			12'd1428 : hue_tab <= 6'd40;
			12'd1429 : hue_tab <= 6'd40;
			12'd1430 : hue_tab <= 6'd40;
			12'd1431 : hue_tab <= 6'd38;
			12'd1432 : hue_tab <= 6'd36;
			12'd1433 : hue_tab <= 6'd35;
			12'd1434 : hue_tab <= 6'd33;
			12'd1435 : hue_tab <= 6'd32;
			12'd1436 : hue_tab <= 6'd31;
			12'd1437 : hue_tab <= 6'd30;
			12'd1438 : hue_tab <= 6'd29;
			12'd1439 : hue_tab <= 6'd28;
			12'd1440 : hue_tab <= 6'd27;
			12'd1441 : hue_tab <= 6'd26;
			12'd1442 : hue_tab <= 6'd25;
			12'd1443 : hue_tab <= 6'd25;
			12'd1444 : hue_tab <= 6'd24;
			12'd1445 : hue_tab <= 6'd23;
			12'd1446 : hue_tab <= 6'd23;
			12'd1447 : hue_tab <= 6'd22;
			12'd1448 : hue_tab <= 6'd22;
			12'd1449 : hue_tab <= 6'd21;
			12'd1450 : hue_tab <= 6'd20;
			12'd1451 : hue_tab <= 6'd20;
			12'd1452 : hue_tab <= 6'd20;
			12'd1453 : hue_tab <= 6'd19;
			12'd1454 : hue_tab <= 6'd19;
			12'd1455 : hue_tab <= 6'd18;
			12'd1456 : hue_tab <= 6'd18;
			12'd1457 : hue_tab <= 6'd17;
			12'd1458 : hue_tab <= 6'd17;
			12'd1459 : hue_tab <= 6'd17;
			12'd1460 : hue_tab <= 6'd16;
			12'd1461 : hue_tab <= 6'd16;
			12'd1462 : hue_tab <= 6'd16;
			12'd1463 : hue_tab <= 6'd16;
			12'd1464 : hue_tab <= 6'd15;
			12'd1465 : hue_tab <= 6'd15;
			12'd1466 : hue_tab <= 6'd15;
			12'd1467 : hue_tab <= 6'd14;
			12'd1468 : hue_tab <= 6'd14;
			12'd1469 : hue_tab <= 6'd14;
			12'd1470 : hue_tab <= 6'd14;
			12'd1471 : hue_tab <= 6'd13;
			12'd1472 : hue_tab <= 6'd0;
			12'd1473 : hue_tab <= 6'd40;
			12'd1474 : hue_tab <= 6'd40;
			12'd1475 : hue_tab <= 6'd40;
			12'd1476 : hue_tab <= 6'd40;
			12'd1477 : hue_tab <= 6'd40;
			12'd1478 : hue_tab <= 6'd40;
			12'd1479 : hue_tab <= 6'd40;
			12'd1480 : hue_tab <= 6'd40;
			12'd1481 : hue_tab <= 6'd40;
			12'd1482 : hue_tab <= 6'd40;
			12'd1483 : hue_tab <= 6'd40;
			12'd1484 : hue_tab <= 6'd40;
			12'd1485 : hue_tab <= 6'd40;
			12'd1486 : hue_tab <= 6'd40;
			12'd1487 : hue_tab <= 6'd40;
			12'd1488 : hue_tab <= 6'd40;
			12'd1489 : hue_tab <= 6'd40;
			12'd1490 : hue_tab <= 6'd40;
			12'd1491 : hue_tab <= 6'd40;
			12'd1492 : hue_tab <= 6'd40;
			12'd1493 : hue_tab <= 6'd40;
			12'd1494 : hue_tab <= 6'd40;
			12'd1495 : hue_tab <= 6'd40;
			12'd1496 : hue_tab <= 6'd38;
			12'd1497 : hue_tab <= 6'd36;
			12'd1498 : hue_tab <= 6'd35;
			12'd1499 : hue_tab <= 6'd34;
			12'd1500 : hue_tab <= 6'd32;
			12'd1501 : hue_tab <= 6'd31;
			12'd1502 : hue_tab <= 6'd30;
			12'd1503 : hue_tab <= 6'd29;
			12'd1504 : hue_tab <= 6'd28;
			12'd1505 : hue_tab <= 6'd27;
			12'd1506 : hue_tab <= 6'd27;
			12'd1507 : hue_tab <= 6'd26;
			12'd1508 : hue_tab <= 6'd25;
			12'd1509 : hue_tab <= 6'd24;
			12'd1510 : hue_tab <= 6'd24;
			12'd1511 : hue_tab <= 6'd23;
			12'd1512 : hue_tab <= 6'd23;
			12'd1513 : hue_tab <= 6'd22;
			12'd1514 : hue_tab <= 6'd21;
			12'd1515 : hue_tab <= 6'd21;
			12'd1516 : hue_tab <= 6'd20;
			12'd1517 : hue_tab <= 6'd20;
			12'd1518 : hue_tab <= 6'd20;
			12'd1519 : hue_tab <= 6'd19;
			12'd1520 : hue_tab <= 6'd19;
			12'd1521 : hue_tab <= 6'd18;
			12'd1522 : hue_tab <= 6'd18;
			12'd1523 : hue_tab <= 6'd18;
			12'd1524 : hue_tab <= 6'd17;
			12'd1525 : hue_tab <= 6'd17;
			12'd1526 : hue_tab <= 6'd17;
			12'd1527 : hue_tab <= 6'd16;
			12'd1528 : hue_tab <= 6'd16;
			12'd1529 : hue_tab <= 6'd16;
			12'd1530 : hue_tab <= 6'd15;
			12'd1531 : hue_tab <= 6'd15;
			12'd1532 : hue_tab <= 6'd15;
			12'd1533 : hue_tab <= 6'd15;
			12'd1534 : hue_tab <= 6'd14;
			12'd1535 : hue_tab <= 6'd14;
			12'd1536 : hue_tab <= 6'd0;
			12'd1537 : hue_tab <= 6'd40;
			12'd1538 : hue_tab <= 6'd40;
			12'd1539 : hue_tab <= 6'd40;
			12'd1540 : hue_tab <= 6'd40;
			12'd1541 : hue_tab <= 6'd40;
			12'd1542 : hue_tab <= 6'd40;
			12'd1543 : hue_tab <= 6'd40;
			12'd1544 : hue_tab <= 6'd40;
			12'd1545 : hue_tab <= 6'd40;
			12'd1546 : hue_tab <= 6'd40;
			12'd1547 : hue_tab <= 6'd40;
			12'd1548 : hue_tab <= 6'd40;
			12'd1549 : hue_tab <= 6'd40;
			12'd1550 : hue_tab <= 6'd40;
			12'd1551 : hue_tab <= 6'd40;
			12'd1552 : hue_tab <= 6'd40;
			12'd1553 : hue_tab <= 6'd40;
			12'd1554 : hue_tab <= 6'd40;
			12'd1555 : hue_tab <= 6'd40;
			12'd1556 : hue_tab <= 6'd40;
			12'd1557 : hue_tab <= 6'd40;
			12'd1558 : hue_tab <= 6'd40;
			12'd1559 : hue_tab <= 6'd40;
			12'd1560 : hue_tab <= 6'd40;
			12'd1561 : hue_tab <= 6'd38;
			12'd1562 : hue_tab <= 6'd36;
			12'd1563 : hue_tab <= 6'd35;
			12'd1564 : hue_tab <= 6'd34;
			12'd1565 : hue_tab <= 6'd33;
			12'd1566 : hue_tab <= 6'd32;
			12'd1567 : hue_tab <= 6'd30;
			12'd1568 : hue_tab <= 6'd30;
			12'd1569 : hue_tab <= 6'd29;
			12'd1570 : hue_tab <= 6'd28;
			12'd1571 : hue_tab <= 6'd27;
			12'd1572 : hue_tab <= 6'd26;
			12'd1573 : hue_tab <= 6'd25;
			12'd1574 : hue_tab <= 6'd25;
			12'd1575 : hue_tab <= 6'd24;
			12'd1576 : hue_tab <= 6'd24;
			12'd1577 : hue_tab <= 6'd23;
			12'd1578 : hue_tab <= 6'd22;
			12'd1579 : hue_tab <= 6'd22;
			12'd1580 : hue_tab <= 6'd21;
			12'd1581 : hue_tab <= 6'd21;
			12'd1582 : hue_tab <= 6'd20;
			12'd1583 : hue_tab <= 6'd20;
			12'd1584 : hue_tab <= 6'd20;
			12'd1585 : hue_tab <= 6'd19;
			12'd1586 : hue_tab <= 6'd19;
			12'd1587 : hue_tab <= 6'd18;
			12'd1588 : hue_tab <= 6'd18;
			12'd1589 : hue_tab <= 6'd18;
			12'd1590 : hue_tab <= 6'd17;
			12'd1591 : hue_tab <= 6'd17;
			12'd1592 : hue_tab <= 6'd17;
			12'd1593 : hue_tab <= 6'd16;
			12'd1594 : hue_tab <= 6'd16;
			12'd1595 : hue_tab <= 6'd16;
			12'd1596 : hue_tab <= 6'd16;
			12'd1597 : hue_tab <= 6'd15;
			12'd1598 : hue_tab <= 6'd15;
			12'd1599 : hue_tab <= 6'd15;
			12'd1600 : hue_tab <= 6'd0;
			12'd1601 : hue_tab <= 6'd40;
			12'd1602 : hue_tab <= 6'd40;
			12'd1603 : hue_tab <= 6'd40;
			12'd1604 : hue_tab <= 6'd40;
			12'd1605 : hue_tab <= 6'd40;
			12'd1606 : hue_tab <= 6'd40;
			12'd1607 : hue_tab <= 6'd40;
			12'd1608 : hue_tab <= 6'd40;
			12'd1609 : hue_tab <= 6'd40;
			12'd1610 : hue_tab <= 6'd40;
			12'd1611 : hue_tab <= 6'd40;
			12'd1612 : hue_tab <= 6'd40;
			12'd1613 : hue_tab <= 6'd40;
			12'd1614 : hue_tab <= 6'd40;
			12'd1615 : hue_tab <= 6'd40;
			12'd1616 : hue_tab <= 6'd40;
			12'd1617 : hue_tab <= 6'd40;
			12'd1618 : hue_tab <= 6'd40;
			12'd1619 : hue_tab <= 6'd40;
			12'd1620 : hue_tab <= 6'd40;
			12'd1621 : hue_tab <= 6'd40;
			12'd1622 : hue_tab <= 6'd40;
			12'd1623 : hue_tab <= 6'd40;
			12'd1624 : hue_tab <= 6'd40;
			12'd1625 : hue_tab <= 6'd40;
			12'd1626 : hue_tab <= 6'd38;
			12'd1627 : hue_tab <= 6'd37;
			12'd1628 : hue_tab <= 6'd35;
			12'd1629 : hue_tab <= 6'd34;
			12'd1630 : hue_tab <= 6'd33;
			12'd1631 : hue_tab <= 6'd32;
			12'd1632 : hue_tab <= 6'd31;
			12'd1633 : hue_tab <= 6'd30;
			12'd1634 : hue_tab <= 6'd29;
			12'd1635 : hue_tab <= 6'd28;
			12'd1636 : hue_tab <= 6'd27;
			12'd1637 : hue_tab <= 6'd27;
			12'd1638 : hue_tab <= 6'd26;
			12'd1639 : hue_tab <= 6'd25;
			12'd1640 : hue_tab <= 6'd25;
			12'd1641 : hue_tab <= 6'd24;
			12'd1642 : hue_tab <= 6'd23;
			12'd1643 : hue_tab <= 6'd23;
			12'd1644 : hue_tab <= 6'd22;
			12'd1645 : hue_tab <= 6'd22;
			12'd1646 : hue_tab <= 6'd21;
			12'd1647 : hue_tab <= 6'd21;
			12'd1648 : hue_tab <= 6'd20;
			12'd1649 : hue_tab <= 6'd20;
			12'd1650 : hue_tab <= 6'd20;
			12'd1651 : hue_tab <= 6'd19;
			12'd1652 : hue_tab <= 6'd19;
			12'd1653 : hue_tab <= 6'd18;
			12'd1654 : hue_tab <= 6'd18;
			12'd1655 : hue_tab <= 6'd18;
			12'd1656 : hue_tab <= 6'd17;
			12'd1657 : hue_tab <= 6'd17;
			12'd1658 : hue_tab <= 6'd17;
			12'd1659 : hue_tab <= 6'd16;
			12'd1660 : hue_tab <= 6'd16;
			12'd1661 : hue_tab <= 6'd16;
			12'd1662 : hue_tab <= 6'd16;
			12'd1663 : hue_tab <= 6'd15;
			12'd1664 : hue_tab <= 6'd0;
			12'd1665 : hue_tab <= 6'd40;
			12'd1666 : hue_tab <= 6'd40;
			12'd1667 : hue_tab <= 6'd40;
			12'd1668 : hue_tab <= 6'd40;
			12'd1669 : hue_tab <= 6'd40;
			12'd1670 : hue_tab <= 6'd40;
			12'd1671 : hue_tab <= 6'd40;
			12'd1672 : hue_tab <= 6'd40;
			12'd1673 : hue_tab <= 6'd40;
			12'd1674 : hue_tab <= 6'd40;
			12'd1675 : hue_tab <= 6'd40;
			12'd1676 : hue_tab <= 6'd40;
			12'd1677 : hue_tab <= 6'd40;
			12'd1678 : hue_tab <= 6'd40;
			12'd1679 : hue_tab <= 6'd40;
			12'd1680 : hue_tab <= 6'd40;
			12'd1681 : hue_tab <= 6'd40;
			12'd1682 : hue_tab <= 6'd40;
			12'd1683 : hue_tab <= 6'd40;
			12'd1684 : hue_tab <= 6'd40;
			12'd1685 : hue_tab <= 6'd40;
			12'd1686 : hue_tab <= 6'd40;
			12'd1687 : hue_tab <= 6'd40;
			12'd1688 : hue_tab <= 6'd40;
			12'd1689 : hue_tab <= 6'd40;
			12'd1690 : hue_tab <= 6'd40;
			12'd1691 : hue_tab <= 6'd38;
			12'd1692 : hue_tab <= 6'd37;
			12'd1693 : hue_tab <= 6'd35;
			12'd1694 : hue_tab <= 6'd34;
			12'd1695 : hue_tab <= 6'd33;
			12'd1696 : hue_tab <= 6'd32;
			12'd1697 : hue_tab <= 6'd31;
			12'd1698 : hue_tab <= 6'd30;
			12'd1699 : hue_tab <= 6'd29;
			12'd1700 : hue_tab <= 6'd28;
			12'd1701 : hue_tab <= 6'd28;
			12'd1702 : hue_tab <= 6'd27;
			12'd1703 : hue_tab <= 6'd26;
			12'd1704 : hue_tab <= 6'd26;
			12'd1705 : hue_tab <= 6'd25;
			12'd1706 : hue_tab <= 6'd24;
			12'd1707 : hue_tab <= 6'd24;
			12'd1708 : hue_tab <= 6'd23;
			12'd1709 : hue_tab <= 6'd23;
			12'd1710 : hue_tab <= 6'd22;
			12'd1711 : hue_tab <= 6'd22;
			12'd1712 : hue_tab <= 6'd21;
			12'd1713 : hue_tab <= 6'd21;
			12'd1714 : hue_tab <= 6'd20;
			12'd1715 : hue_tab <= 6'd20;
			12'd1716 : hue_tab <= 6'd20;
			12'd1717 : hue_tab <= 6'd19;
			12'd1718 : hue_tab <= 6'd19;
			12'd1719 : hue_tab <= 6'd18;
			12'd1720 : hue_tab <= 6'd18;
			12'd1721 : hue_tab <= 6'd18;
			12'd1722 : hue_tab <= 6'd17;
			12'd1723 : hue_tab <= 6'd17;
			12'd1724 : hue_tab <= 6'd17;
			12'd1725 : hue_tab <= 6'd17;
			12'd1726 : hue_tab <= 6'd16;
			12'd1727 : hue_tab <= 6'd16;
			12'd1728 : hue_tab <= 6'd0;
			12'd1729 : hue_tab <= 6'd40;
			12'd1730 : hue_tab <= 6'd40;
			12'd1731 : hue_tab <= 6'd40;
			12'd1732 : hue_tab <= 6'd40;
			12'd1733 : hue_tab <= 6'd40;
			12'd1734 : hue_tab <= 6'd40;
			12'd1735 : hue_tab <= 6'd40;
			12'd1736 : hue_tab <= 6'd40;
			12'd1737 : hue_tab <= 6'd40;
			12'd1738 : hue_tab <= 6'd40;
			12'd1739 : hue_tab <= 6'd40;
			12'd1740 : hue_tab <= 6'd40;
			12'd1741 : hue_tab <= 6'd40;
			12'd1742 : hue_tab <= 6'd40;
			12'd1743 : hue_tab <= 6'd40;
			12'd1744 : hue_tab <= 6'd40;
			12'd1745 : hue_tab <= 6'd40;
			12'd1746 : hue_tab <= 6'd40;
			12'd1747 : hue_tab <= 6'd40;
			12'd1748 : hue_tab <= 6'd40;
			12'd1749 : hue_tab <= 6'd40;
			12'd1750 : hue_tab <= 6'd40;
			12'd1751 : hue_tab <= 6'd40;
			12'd1752 : hue_tab <= 6'd40;
			12'd1753 : hue_tab <= 6'd40;
			12'd1754 : hue_tab <= 6'd40;
			12'd1755 : hue_tab <= 6'd40;
			12'd1756 : hue_tab <= 6'd38;
			12'd1757 : hue_tab <= 6'd37;
			12'd1758 : hue_tab <= 6'd36;
			12'd1759 : hue_tab <= 6'd34;
			12'd1760 : hue_tab <= 6'd33;
			12'd1761 : hue_tab <= 6'd32;
			12'd1762 : hue_tab <= 6'd31;
			12'd1763 : hue_tab <= 6'd30;
			12'd1764 : hue_tab <= 6'd30;
			12'd1765 : hue_tab <= 6'd29;
			12'd1766 : hue_tab <= 6'd28;
			12'd1767 : hue_tab <= 6'd27;
			12'd1768 : hue_tab <= 6'd27;
			12'd1769 : hue_tab <= 6'd26;
			12'd1770 : hue_tab <= 6'd25;
			12'd1771 : hue_tab <= 6'd25;
			12'd1772 : hue_tab <= 6'd24;
			12'd1773 : hue_tab <= 6'd24;
			12'd1774 : hue_tab <= 6'd23;
			12'd1775 : hue_tab <= 6'd22;
			12'd1776 : hue_tab <= 6'd22;
			12'd1777 : hue_tab <= 6'd22;
			12'd1778 : hue_tab <= 6'd21;
			12'd1779 : hue_tab <= 6'd21;
			12'd1780 : hue_tab <= 6'd20;
			12'd1781 : hue_tab <= 6'd20;
			12'd1782 : hue_tab <= 6'd20;
			12'd1783 : hue_tab <= 6'd19;
			12'd1784 : hue_tab <= 6'd19;
			12'd1785 : hue_tab <= 6'd18;
			12'd1786 : hue_tab <= 6'd18;
			12'd1787 : hue_tab <= 6'd18;
			12'd1788 : hue_tab <= 6'd18;
			12'd1789 : hue_tab <= 6'd17;
			12'd1790 : hue_tab <= 6'd17;
			12'd1791 : hue_tab <= 6'd17;
			12'd1792 : hue_tab <= 6'd0;
			12'd1793 : hue_tab <= 6'd40;
			12'd1794 : hue_tab <= 6'd40;
			12'd1795 : hue_tab <= 6'd40;
			12'd1796 : hue_tab <= 6'd40;
			12'd1797 : hue_tab <= 6'd40;
			12'd1798 : hue_tab <= 6'd40;
			12'd1799 : hue_tab <= 6'd40;
			12'd1800 : hue_tab <= 6'd40;
			12'd1801 : hue_tab <= 6'd40;
			12'd1802 : hue_tab <= 6'd40;
			12'd1803 : hue_tab <= 6'd40;
			12'd1804 : hue_tab <= 6'd40;
			12'd1805 : hue_tab <= 6'd40;
			12'd1806 : hue_tab <= 6'd40;
			12'd1807 : hue_tab <= 6'd40;
			12'd1808 : hue_tab <= 6'd40;
			12'd1809 : hue_tab <= 6'd40;
			12'd1810 : hue_tab <= 6'd40;
			12'd1811 : hue_tab <= 6'd40;
			12'd1812 : hue_tab <= 6'd40;
			12'd1813 : hue_tab <= 6'd40;
			12'd1814 : hue_tab <= 6'd40;
			12'd1815 : hue_tab <= 6'd40;
			12'd1816 : hue_tab <= 6'd40;
			12'd1817 : hue_tab <= 6'd40;
			12'd1818 : hue_tab <= 6'd40;
			12'd1819 : hue_tab <= 6'd40;
			12'd1820 : hue_tab <= 6'd40;
			12'd1821 : hue_tab <= 6'd38;
			12'd1822 : hue_tab <= 6'd37;
			12'd1823 : hue_tab <= 6'd36;
			12'd1824 : hue_tab <= 6'd35;
			12'd1825 : hue_tab <= 6'd33;
			12'd1826 : hue_tab <= 6'd32;
			12'd1827 : hue_tab <= 6'd32;
			12'd1828 : hue_tab <= 6'd31;
			12'd1829 : hue_tab <= 6'd30;
			12'd1830 : hue_tab <= 6'd29;
			12'd1831 : hue_tab <= 6'd28;
			12'd1832 : hue_tab <= 6'd28;
			12'd1833 : hue_tab <= 6'd27;
			12'd1834 : hue_tab <= 6'd26;
			12'd1835 : hue_tab <= 6'd26;
			12'd1836 : hue_tab <= 6'd25;
			12'd1837 : hue_tab <= 6'd24;
			12'd1838 : hue_tab <= 6'd24;
			12'd1839 : hue_tab <= 6'd23;
			12'd1840 : hue_tab <= 6'd23;
			12'd1841 : hue_tab <= 6'd22;
			12'd1842 : hue_tab <= 6'd22;
			12'd1843 : hue_tab <= 6'd21;
			12'd1844 : hue_tab <= 6'd21;
			12'd1845 : hue_tab <= 6'd21;
			12'd1846 : hue_tab <= 6'd20;
			12'd1847 : hue_tab <= 6'd20;
			12'd1848 : hue_tab <= 6'd20;
			12'd1849 : hue_tab <= 6'd19;
			12'd1850 : hue_tab <= 6'd19;
			12'd1851 : hue_tab <= 6'd18;
			12'd1852 : hue_tab <= 6'd18;
			12'd1853 : hue_tab <= 6'd18;
			12'd1854 : hue_tab <= 6'd18;
			12'd1855 : hue_tab <= 6'd17;
			12'd1856 : hue_tab <= 6'd0;
			12'd1857 : hue_tab <= 6'd40;
			12'd1858 : hue_tab <= 6'd40;
			12'd1859 : hue_tab <= 6'd40;
			12'd1860 : hue_tab <= 6'd40;
			12'd1861 : hue_tab <= 6'd40;
			12'd1862 : hue_tab <= 6'd40;
			12'd1863 : hue_tab <= 6'd40;
			12'd1864 : hue_tab <= 6'd40;
			12'd1865 : hue_tab <= 6'd40;
			12'd1866 : hue_tab <= 6'd40;
			12'd1867 : hue_tab <= 6'd40;
			12'd1868 : hue_tab <= 6'd40;
			12'd1869 : hue_tab <= 6'd40;
			12'd1870 : hue_tab <= 6'd40;
			12'd1871 : hue_tab <= 6'd40;
			12'd1872 : hue_tab <= 6'd40;
			12'd1873 : hue_tab <= 6'd40;
			12'd1874 : hue_tab <= 6'd40;
			12'd1875 : hue_tab <= 6'd40;
			12'd1876 : hue_tab <= 6'd40;
			12'd1877 : hue_tab <= 6'd40;
			12'd1878 : hue_tab <= 6'd40;
			12'd1879 : hue_tab <= 6'd40;
			12'd1880 : hue_tab <= 6'd40;
			12'd1881 : hue_tab <= 6'd40;
			12'd1882 : hue_tab <= 6'd40;
			12'd1883 : hue_tab <= 6'd40;
			12'd1884 : hue_tab <= 6'd40;
			12'd1885 : hue_tab <= 6'd40;
			12'd1886 : hue_tab <= 6'd38;
			12'd1887 : hue_tab <= 6'd37;
			12'd1888 : hue_tab <= 6'd36;
			12'd1889 : hue_tab <= 6'd35;
			12'd1890 : hue_tab <= 6'd34;
			12'd1891 : hue_tab <= 6'd33;
			12'd1892 : hue_tab <= 6'd32;
			12'd1893 : hue_tab <= 6'd31;
			12'd1894 : hue_tab <= 6'd30;
			12'd1895 : hue_tab <= 6'd29;
			12'd1896 : hue_tab <= 6'd29;
			12'd1897 : hue_tab <= 6'd28;
			12'd1898 : hue_tab <= 6'd27;
			12'd1899 : hue_tab <= 6'd26;
			12'd1900 : hue_tab <= 6'd26;
			12'd1901 : hue_tab <= 6'd25;
			12'd1902 : hue_tab <= 6'd25;
			12'd1903 : hue_tab <= 6'd24;
			12'd1904 : hue_tab <= 6'd24;
			12'd1905 : hue_tab <= 6'd23;
			12'd1906 : hue_tab <= 6'd23;
			12'd1907 : hue_tab <= 6'd22;
			12'd1908 : hue_tab <= 6'd22;
			12'd1909 : hue_tab <= 6'd21;
			12'd1910 : hue_tab <= 6'd21;
			12'd1911 : hue_tab <= 6'd21;
			12'd1912 : hue_tab <= 6'd20;
			12'd1913 : hue_tab <= 6'd20;
			12'd1914 : hue_tab <= 6'd20;
			12'd1915 : hue_tab <= 6'd19;
			12'd1916 : hue_tab <= 6'd19;
			12'd1917 : hue_tab <= 6'd19;
			12'd1918 : hue_tab <= 6'd18;
			12'd1919 : hue_tab <= 6'd18;
			12'd1920 : hue_tab <= 6'd0;
			12'd1921 : hue_tab <= 6'd40;
			12'd1922 : hue_tab <= 6'd40;
			12'd1923 : hue_tab <= 6'd40;
			12'd1924 : hue_tab <= 6'd40;
			12'd1925 : hue_tab <= 6'd40;
			12'd1926 : hue_tab <= 6'd40;
			12'd1927 : hue_tab <= 6'd40;
			12'd1928 : hue_tab <= 6'd40;
			12'd1929 : hue_tab <= 6'd40;
			12'd1930 : hue_tab <= 6'd40;
			12'd1931 : hue_tab <= 6'd40;
			12'd1932 : hue_tab <= 6'd40;
			12'd1933 : hue_tab <= 6'd40;
			12'd1934 : hue_tab <= 6'd40;
			12'd1935 : hue_tab <= 6'd40;
			12'd1936 : hue_tab <= 6'd40;
			12'd1937 : hue_tab <= 6'd40;
			12'd1938 : hue_tab <= 6'd40;
			12'd1939 : hue_tab <= 6'd40;
			12'd1940 : hue_tab <= 6'd40;
			12'd1941 : hue_tab <= 6'd40;
			12'd1942 : hue_tab <= 6'd40;
			12'd1943 : hue_tab <= 6'd40;
			12'd1944 : hue_tab <= 6'd40;
			12'd1945 : hue_tab <= 6'd40;
			12'd1946 : hue_tab <= 6'd40;
			12'd1947 : hue_tab <= 6'd40;
			12'd1948 : hue_tab <= 6'd40;
			12'd1949 : hue_tab <= 6'd40;
			12'd1950 : hue_tab <= 6'd40;
			12'd1951 : hue_tab <= 6'd38;
			12'd1952 : hue_tab <= 6'd37;
			12'd1953 : hue_tab <= 6'd36;
			12'd1954 : hue_tab <= 6'd35;
			12'd1955 : hue_tab <= 6'd34;
			12'd1956 : hue_tab <= 6'd33;
			12'd1957 : hue_tab <= 6'd32;
			12'd1958 : hue_tab <= 6'd31;
			12'd1959 : hue_tab <= 6'd30;
			12'd1960 : hue_tab <= 6'd30;
			12'd1961 : hue_tab <= 6'd29;
			12'd1962 : hue_tab <= 6'd28;
			12'd1963 : hue_tab <= 6'd27;
			12'd1964 : hue_tab <= 6'd27;
			12'd1965 : hue_tab <= 6'd26;
			12'd1966 : hue_tab <= 6'd26;
			12'd1967 : hue_tab <= 6'd25;
			12'd1968 : hue_tab <= 6'd25;
			12'd1969 : hue_tab <= 6'd24;
			12'd1970 : hue_tab <= 6'd24;
			12'd1971 : hue_tab <= 6'd23;
			12'd1972 : hue_tab <= 6'd23;
			12'd1973 : hue_tab <= 6'd22;
			12'd1974 : hue_tab <= 6'd22;
			12'd1975 : hue_tab <= 6'd21;
			12'd1976 : hue_tab <= 6'd21;
			12'd1977 : hue_tab <= 6'd21;
			12'd1978 : hue_tab <= 6'd20;
			12'd1979 : hue_tab <= 6'd20;
			12'd1980 : hue_tab <= 6'd20;
			12'd1981 : hue_tab <= 6'd19;
			12'd1982 : hue_tab <= 6'd19;
			12'd1983 : hue_tab <= 6'd19;
			12'd1984 : hue_tab <= 6'd0;
			12'd1985 : hue_tab <= 6'd40;
			12'd1986 : hue_tab <= 6'd40;
			12'd1987 : hue_tab <= 6'd40;
			12'd1988 : hue_tab <= 6'd40;
			12'd1989 : hue_tab <= 6'd40;
			12'd1990 : hue_tab <= 6'd40;
			12'd1991 : hue_tab <= 6'd40;
			12'd1992 : hue_tab <= 6'd40;
			12'd1993 : hue_tab <= 6'd40;
			12'd1994 : hue_tab <= 6'd40;
			12'd1995 : hue_tab <= 6'd40;
			12'd1996 : hue_tab <= 6'd40;
			12'd1997 : hue_tab <= 6'd40;
			12'd1998 : hue_tab <= 6'd40;
			12'd1999 : hue_tab <= 6'd40;
			12'd2000 : hue_tab <= 6'd40;
			12'd2001 : hue_tab <= 6'd40;
			12'd2002 : hue_tab <= 6'd40;
			12'd2003 : hue_tab <= 6'd40;
			12'd2004 : hue_tab <= 6'd40;
			12'd2005 : hue_tab <= 6'd40;
			12'd2006 : hue_tab <= 6'd40;
			12'd2007 : hue_tab <= 6'd40;
			12'd2008 : hue_tab <= 6'd40;
			12'd2009 : hue_tab <= 6'd40;
			12'd2010 : hue_tab <= 6'd40;
			12'd2011 : hue_tab <= 6'd40;
			12'd2012 : hue_tab <= 6'd40;
			12'd2013 : hue_tab <= 6'd40;
			12'd2014 : hue_tab <= 6'd40;
			12'd2015 : hue_tab <= 6'd40;
			12'd2016 : hue_tab <= 6'd38;
			12'd2017 : hue_tab <= 6'd37;
			12'd2018 : hue_tab <= 6'd36;
			12'd2019 : hue_tab <= 6'd35;
			12'd2020 : hue_tab <= 6'd34;
			12'd2021 : hue_tab <= 6'd33;
			12'd2022 : hue_tab <= 6'd32;
			12'd2023 : hue_tab <= 6'd31;
			12'd2024 : hue_tab <= 6'd31;
			12'd2025 : hue_tab <= 6'd30;
			12'd2026 : hue_tab <= 6'd29;
			12'd2027 : hue_tab <= 6'd28;
			12'd2028 : hue_tab <= 6'd28;
			12'd2029 : hue_tab <= 6'd27;
			12'd2030 : hue_tab <= 6'd26;
			12'd2031 : hue_tab <= 6'd26;
			12'd2032 : hue_tab <= 6'd25;
			12'd2033 : hue_tab <= 6'd25;
			12'd2034 : hue_tab <= 6'd24;
			12'd2035 : hue_tab <= 6'd24;
			12'd2036 : hue_tab <= 6'd23;
			12'd2037 : hue_tab <= 6'd23;
			12'd2038 : hue_tab <= 6'd22;
			12'd2039 : hue_tab <= 6'd22;
			12'd2040 : hue_tab <= 6'd22;
			12'd2041 : hue_tab <= 6'd21;
			12'd2042 : hue_tab <= 6'd21;
			12'd2043 : hue_tab <= 6'd21;
			12'd2044 : hue_tab <= 6'd20;
			12'd2045 : hue_tab <= 6'd20;
			12'd2046 : hue_tab <= 6'd20;
			12'd2047 : hue_tab <= 6'd19;
			12'd2048 : hue_tab <= 6'd0;
			12'd2049 : hue_tab <= 6'd40;
			12'd2050 : hue_tab <= 6'd40;
			12'd2051 : hue_tab <= 6'd40;
			12'd2052 : hue_tab <= 6'd40;
			12'd2053 : hue_tab <= 6'd40;
			12'd2054 : hue_tab <= 6'd40;
			12'd2055 : hue_tab <= 6'd40;
			12'd2056 : hue_tab <= 6'd40;
			12'd2057 : hue_tab <= 6'd40;
			12'd2058 : hue_tab <= 6'd40;
			12'd2059 : hue_tab <= 6'd40;
			12'd2060 : hue_tab <= 6'd40;
			12'd2061 : hue_tab <= 6'd40;
			12'd2062 : hue_tab <= 6'd40;
			12'd2063 : hue_tab <= 6'd40;
			12'd2064 : hue_tab <= 6'd40;
			12'd2065 : hue_tab <= 6'd40;
			12'd2066 : hue_tab <= 6'd40;
			12'd2067 : hue_tab <= 6'd40;
			12'd2068 : hue_tab <= 6'd40;
			12'd2069 : hue_tab <= 6'd40;
			12'd2070 : hue_tab <= 6'd40;
			12'd2071 : hue_tab <= 6'd40;
			12'd2072 : hue_tab <= 6'd40;
			12'd2073 : hue_tab <= 6'd40;
			12'd2074 : hue_tab <= 6'd40;
			12'd2075 : hue_tab <= 6'd40;
			12'd2076 : hue_tab <= 6'd40;
			12'd2077 : hue_tab <= 6'd40;
			12'd2078 : hue_tab <= 6'd40;
			12'd2079 : hue_tab <= 6'd40;
			12'd2080 : hue_tab <= 6'd40;
			12'd2081 : hue_tab <= 6'd38;
			12'd2082 : hue_tab <= 6'd37;
			12'd2083 : hue_tab <= 6'd36;
			12'd2084 : hue_tab <= 6'd35;
			12'd2085 : hue_tab <= 6'd34;
			12'd2086 : hue_tab <= 6'd33;
			12'd2087 : hue_tab <= 6'd32;
			12'd2088 : hue_tab <= 6'd32;
			12'd2089 : hue_tab <= 6'd31;
			12'd2090 : hue_tab <= 6'd30;
			12'd2091 : hue_tab <= 6'd29;
			12'd2092 : hue_tab <= 6'd29;
			12'd2093 : hue_tab <= 6'd28;
			12'd2094 : hue_tab <= 6'd27;
			12'd2095 : hue_tab <= 6'd27;
			12'd2096 : hue_tab <= 6'd26;
			12'd2097 : hue_tab <= 6'd26;
			12'd2098 : hue_tab <= 6'd25;
			12'd2099 : hue_tab <= 6'd25;
			12'd2100 : hue_tab <= 6'd24;
			12'd2101 : hue_tab <= 6'd24;
			12'd2102 : hue_tab <= 6'd23;
			12'd2103 : hue_tab <= 6'd23;
			12'd2104 : hue_tab <= 6'd22;
			12'd2105 : hue_tab <= 6'd22;
			12'd2106 : hue_tab <= 6'd22;
			12'd2107 : hue_tab <= 6'd21;
			12'd2108 : hue_tab <= 6'd21;
			12'd2109 : hue_tab <= 6'd20;
			12'd2110 : hue_tab <= 6'd20;
			12'd2111 : hue_tab <= 6'd20;
			12'd2112 : hue_tab <= 6'd0;
			12'd2113 : hue_tab <= 6'd40;
			12'd2114 : hue_tab <= 6'd40;
			12'd2115 : hue_tab <= 6'd40;
			12'd2116 : hue_tab <= 6'd40;
			12'd2117 : hue_tab <= 6'd40;
			12'd2118 : hue_tab <= 6'd40;
			12'd2119 : hue_tab <= 6'd40;
			12'd2120 : hue_tab <= 6'd40;
			12'd2121 : hue_tab <= 6'd40;
			12'd2122 : hue_tab <= 6'd40;
			12'd2123 : hue_tab <= 6'd40;
			12'd2124 : hue_tab <= 6'd40;
			12'd2125 : hue_tab <= 6'd40;
			12'd2126 : hue_tab <= 6'd40;
			12'd2127 : hue_tab <= 6'd40;
			12'd2128 : hue_tab <= 6'd40;
			12'd2129 : hue_tab <= 6'd40;
			12'd2130 : hue_tab <= 6'd40;
			12'd2131 : hue_tab <= 6'd40;
			12'd2132 : hue_tab <= 6'd40;
			12'd2133 : hue_tab <= 6'd40;
			12'd2134 : hue_tab <= 6'd40;
			12'd2135 : hue_tab <= 6'd40;
			12'd2136 : hue_tab <= 6'd40;
			12'd2137 : hue_tab <= 6'd40;
			12'd2138 : hue_tab <= 6'd40;
			12'd2139 : hue_tab <= 6'd40;
			12'd2140 : hue_tab <= 6'd40;
			12'd2141 : hue_tab <= 6'd40;
			12'd2142 : hue_tab <= 6'd40;
			12'd2143 : hue_tab <= 6'd40;
			12'd2144 : hue_tab <= 6'd40;
			12'd2145 : hue_tab <= 6'd40;
			12'd2146 : hue_tab <= 6'd38;
			12'd2147 : hue_tab <= 6'd37;
			12'd2148 : hue_tab <= 6'd36;
			12'd2149 : hue_tab <= 6'd35;
			12'd2150 : hue_tab <= 6'd34;
			12'd2151 : hue_tab <= 6'd33;
			12'd2152 : hue_tab <= 6'd33;
			12'd2153 : hue_tab <= 6'd32;
			12'd2154 : hue_tab <= 6'd31;
			12'd2155 : hue_tab <= 6'd30;
			12'd2156 : hue_tab <= 6'd30;
			12'd2157 : hue_tab <= 6'd29;
			12'd2158 : hue_tab <= 6'd28;
			12'd2159 : hue_tab <= 6'd28;
			12'd2160 : hue_tab <= 6'd27;
			12'd2161 : hue_tab <= 6'd26;
			12'd2162 : hue_tab <= 6'd26;
			12'd2163 : hue_tab <= 6'd25;
			12'd2164 : hue_tab <= 6'd25;
			12'd2165 : hue_tab <= 6'd24;
			12'd2166 : hue_tab <= 6'd24;
			12'd2167 : hue_tab <= 6'd24;
			12'd2168 : hue_tab <= 6'd23;
			12'd2169 : hue_tab <= 6'd23;
			12'd2170 : hue_tab <= 6'd22;
			12'd2171 : hue_tab <= 6'd22;
			12'd2172 : hue_tab <= 6'd22;
			12'd2173 : hue_tab <= 6'd21;
			12'd2174 : hue_tab <= 6'd21;
			12'd2175 : hue_tab <= 6'd20;
			12'd2176 : hue_tab <= 6'd0;
			12'd2177 : hue_tab <= 6'd40;
			12'd2178 : hue_tab <= 6'd40;
			12'd2179 : hue_tab <= 6'd40;
			12'd2180 : hue_tab <= 6'd40;
			12'd2181 : hue_tab <= 6'd40;
			12'd2182 : hue_tab <= 6'd40;
			12'd2183 : hue_tab <= 6'd40;
			12'd2184 : hue_tab <= 6'd40;
			12'd2185 : hue_tab <= 6'd40;
			12'd2186 : hue_tab <= 6'd40;
			12'd2187 : hue_tab <= 6'd40;
			12'd2188 : hue_tab <= 6'd40;
			12'd2189 : hue_tab <= 6'd40;
			12'd2190 : hue_tab <= 6'd40;
			12'd2191 : hue_tab <= 6'd40;
			12'd2192 : hue_tab <= 6'd40;
			12'd2193 : hue_tab <= 6'd40;
			12'd2194 : hue_tab <= 6'd40;
			12'd2195 : hue_tab <= 6'd40;
			12'd2196 : hue_tab <= 6'd40;
			12'd2197 : hue_tab <= 6'd40;
			12'd2198 : hue_tab <= 6'd40;
			12'd2199 : hue_tab <= 6'd40;
			12'd2200 : hue_tab <= 6'd40;
			12'd2201 : hue_tab <= 6'd40;
			12'd2202 : hue_tab <= 6'd40;
			12'd2203 : hue_tab <= 6'd40;
			12'd2204 : hue_tab <= 6'd40;
			12'd2205 : hue_tab <= 6'd40;
			12'd2206 : hue_tab <= 6'd40;
			12'd2207 : hue_tab <= 6'd40;
			12'd2208 : hue_tab <= 6'd40;
			12'd2209 : hue_tab <= 6'd40;
			12'd2210 : hue_tab <= 6'd40;
			12'd2211 : hue_tab <= 6'd38;
			12'd2212 : hue_tab <= 6'd37;
			12'd2213 : hue_tab <= 6'd36;
			12'd2214 : hue_tab <= 6'd35;
			12'd2215 : hue_tab <= 6'd34;
			12'd2216 : hue_tab <= 6'd34;
			12'd2217 : hue_tab <= 6'd33;
			12'd2218 : hue_tab <= 6'd32;
			12'd2219 : hue_tab <= 6'd31;
			12'd2220 : hue_tab <= 6'd30;
			12'd2221 : hue_tab <= 6'd30;
			12'd2222 : hue_tab <= 6'd29;
			12'd2223 : hue_tab <= 6'd28;
			12'd2224 : hue_tab <= 6'd28;
			12'd2225 : hue_tab <= 6'd27;
			12'd2226 : hue_tab <= 6'd27;
			12'd2227 : hue_tab <= 6'd26;
			12'd2228 : hue_tab <= 6'd26;
			12'd2229 : hue_tab <= 6'd25;
			12'd2230 : hue_tab <= 6'd25;
			12'd2231 : hue_tab <= 6'd24;
			12'd2232 : hue_tab <= 6'd24;
			12'd2233 : hue_tab <= 6'd23;
			12'd2234 : hue_tab <= 6'd23;
			12'd2235 : hue_tab <= 6'd23;
			12'd2236 : hue_tab <= 6'd22;
			12'd2237 : hue_tab <= 6'd22;
			12'd2238 : hue_tab <= 6'd21;
			12'd2239 : hue_tab <= 6'd21;
			12'd2240 : hue_tab <= 6'd0;
			12'd2241 : hue_tab <= 6'd40;
			12'd2242 : hue_tab <= 6'd40;
			12'd2243 : hue_tab <= 6'd40;
			12'd2244 : hue_tab <= 6'd40;
			12'd2245 : hue_tab <= 6'd40;
			12'd2246 : hue_tab <= 6'd40;
			12'd2247 : hue_tab <= 6'd40;
			12'd2248 : hue_tab <= 6'd40;
			12'd2249 : hue_tab <= 6'd40;
			12'd2250 : hue_tab <= 6'd40;
			12'd2251 : hue_tab <= 6'd40;
			12'd2252 : hue_tab <= 6'd40;
			12'd2253 : hue_tab <= 6'd40;
			12'd2254 : hue_tab <= 6'd40;
			12'd2255 : hue_tab <= 6'd40;
			12'd2256 : hue_tab <= 6'd40;
			12'd2257 : hue_tab <= 6'd40;
			12'd2258 : hue_tab <= 6'd40;
			12'd2259 : hue_tab <= 6'd40;
			12'd2260 : hue_tab <= 6'd40;
			12'd2261 : hue_tab <= 6'd40;
			12'd2262 : hue_tab <= 6'd40;
			12'd2263 : hue_tab <= 6'd40;
			12'd2264 : hue_tab <= 6'd40;
			12'd2265 : hue_tab <= 6'd40;
			12'd2266 : hue_tab <= 6'd40;
			12'd2267 : hue_tab <= 6'd40;
			12'd2268 : hue_tab <= 6'd40;
			12'd2269 : hue_tab <= 6'd40;
			12'd2270 : hue_tab <= 6'd40;
			12'd2271 : hue_tab <= 6'd40;
			12'd2272 : hue_tab <= 6'd40;
			12'd2273 : hue_tab <= 6'd40;
			12'd2274 : hue_tab <= 6'd40;
			12'd2275 : hue_tab <= 6'd40;
			12'd2276 : hue_tab <= 6'd38;
			12'd2277 : hue_tab <= 6'd37;
			12'd2278 : hue_tab <= 6'd36;
			12'd2279 : hue_tab <= 6'd35;
			12'd2280 : hue_tab <= 6'd35;
			12'd2281 : hue_tab <= 6'd34;
			12'd2282 : hue_tab <= 6'd33;
			12'd2283 : hue_tab <= 6'd32;
			12'd2284 : hue_tab <= 6'd31;
			12'd2285 : hue_tab <= 6'd31;
			12'd2286 : hue_tab <= 6'd30;
			12'd2287 : hue_tab <= 6'd29;
			12'd2288 : hue_tab <= 6'd29;
			12'd2289 : hue_tab <= 6'd28;
			12'd2290 : hue_tab <= 6'd28;
			12'd2291 : hue_tab <= 6'd27;
			12'd2292 : hue_tab <= 6'd26;
			12'd2293 : hue_tab <= 6'd26;
			12'd2294 : hue_tab <= 6'd25;
			12'd2295 : hue_tab <= 6'd25;
			12'd2296 : hue_tab <= 6'd25;
			12'd2297 : hue_tab <= 6'd24;
			12'd2298 : hue_tab <= 6'd24;
			12'd2299 : hue_tab <= 6'd23;
			12'd2300 : hue_tab <= 6'd23;
			12'd2301 : hue_tab <= 6'd22;
			12'd2302 : hue_tab <= 6'd22;
			12'd2303 : hue_tab <= 6'd22;
			12'd2304 : hue_tab <= 6'd0;
			12'd2305 : hue_tab <= 6'd40;
			12'd2306 : hue_tab <= 6'd40;
			12'd2307 : hue_tab <= 6'd40;
			12'd2308 : hue_tab <= 6'd40;
			12'd2309 : hue_tab <= 6'd40;
			12'd2310 : hue_tab <= 6'd40;
			12'd2311 : hue_tab <= 6'd40;
			12'd2312 : hue_tab <= 6'd40;
			12'd2313 : hue_tab <= 6'd40;
			12'd2314 : hue_tab <= 6'd40;
			12'd2315 : hue_tab <= 6'd40;
			12'd2316 : hue_tab <= 6'd40;
			12'd2317 : hue_tab <= 6'd40;
			12'd2318 : hue_tab <= 6'd40;
			12'd2319 : hue_tab <= 6'd40;
			12'd2320 : hue_tab <= 6'd40;
			12'd2321 : hue_tab <= 6'd40;
			12'd2322 : hue_tab <= 6'd40;
			12'd2323 : hue_tab <= 6'd40;
			12'd2324 : hue_tab <= 6'd40;
			12'd2325 : hue_tab <= 6'd40;
			12'd2326 : hue_tab <= 6'd40;
			12'd2327 : hue_tab <= 6'd40;
			12'd2328 : hue_tab <= 6'd40;
			12'd2329 : hue_tab <= 6'd40;
			12'd2330 : hue_tab <= 6'd40;
			12'd2331 : hue_tab <= 6'd40;
			12'd2332 : hue_tab <= 6'd40;
			12'd2333 : hue_tab <= 6'd40;
			12'd2334 : hue_tab <= 6'd40;
			12'd2335 : hue_tab <= 6'd40;
			12'd2336 : hue_tab <= 6'd40;
			12'd2337 : hue_tab <= 6'd40;
			12'd2338 : hue_tab <= 6'd40;
			12'd2339 : hue_tab <= 6'd40;
			12'd2340 : hue_tab <= 6'd40;
			12'd2341 : hue_tab <= 6'd38;
			12'd2342 : hue_tab <= 6'd37;
			12'd2343 : hue_tab <= 6'd36;
			12'd2344 : hue_tab <= 6'd36;
			12'd2345 : hue_tab <= 6'd35;
			12'd2346 : hue_tab <= 6'd34;
			12'd2347 : hue_tab <= 6'd33;
			12'd2348 : hue_tab <= 6'd32;
			12'd2349 : hue_tab <= 6'd32;
			12'd2350 : hue_tab <= 6'd31;
			12'd2351 : hue_tab <= 6'd30;
			12'd2352 : hue_tab <= 6'd30;
			12'd2353 : hue_tab <= 6'd29;
			12'd2354 : hue_tab <= 6'd28;
			12'd2355 : hue_tab <= 6'd28;
			12'd2356 : hue_tab <= 6'd27;
			12'd2357 : hue_tab <= 6'd27;
			12'd2358 : hue_tab <= 6'd26;
			12'd2359 : hue_tab <= 6'd26;
			12'd2360 : hue_tab <= 6'd25;
			12'd2361 : hue_tab <= 6'd25;
			12'd2362 : hue_tab <= 6'd24;
			12'd2363 : hue_tab <= 6'd24;
			12'd2364 : hue_tab <= 6'd24;
			12'd2365 : hue_tab <= 6'd23;
			12'd2366 : hue_tab <= 6'd23;
			12'd2367 : hue_tab <= 6'd22;
			12'd2368 : hue_tab <= 6'd0;
			12'd2369 : hue_tab <= 6'd40;
			12'd2370 : hue_tab <= 6'd40;
			12'd2371 : hue_tab <= 6'd40;
			12'd2372 : hue_tab <= 6'd40;
			12'd2373 : hue_tab <= 6'd40;
			12'd2374 : hue_tab <= 6'd40;
			12'd2375 : hue_tab <= 6'd40;
			12'd2376 : hue_tab <= 6'd40;
			12'd2377 : hue_tab <= 6'd40;
			12'd2378 : hue_tab <= 6'd40;
			12'd2379 : hue_tab <= 6'd40;
			12'd2380 : hue_tab <= 6'd40;
			12'd2381 : hue_tab <= 6'd40;
			12'd2382 : hue_tab <= 6'd40;
			12'd2383 : hue_tab <= 6'd40;
			12'd2384 : hue_tab <= 6'd40;
			12'd2385 : hue_tab <= 6'd40;
			12'd2386 : hue_tab <= 6'd40;
			12'd2387 : hue_tab <= 6'd40;
			12'd2388 : hue_tab <= 6'd40;
			12'd2389 : hue_tab <= 6'd40;
			12'd2390 : hue_tab <= 6'd40;
			12'd2391 : hue_tab <= 6'd40;
			12'd2392 : hue_tab <= 6'd40;
			12'd2393 : hue_tab <= 6'd40;
			12'd2394 : hue_tab <= 6'd40;
			12'd2395 : hue_tab <= 6'd40;
			12'd2396 : hue_tab <= 6'd40;
			12'd2397 : hue_tab <= 6'd40;
			12'd2398 : hue_tab <= 6'd40;
			12'd2399 : hue_tab <= 6'd40;
			12'd2400 : hue_tab <= 6'd40;
			12'd2401 : hue_tab <= 6'd40;
			12'd2402 : hue_tab <= 6'd40;
			12'd2403 : hue_tab <= 6'd40;
			12'd2404 : hue_tab <= 6'd40;
			12'd2405 : hue_tab <= 6'd40;
			12'd2406 : hue_tab <= 6'd38;
			12'd2407 : hue_tab <= 6'd37;
			12'd2408 : hue_tab <= 6'd37;
			12'd2409 : hue_tab <= 6'd36;
			12'd2410 : hue_tab <= 6'd35;
			12'd2411 : hue_tab <= 6'd34;
			12'd2412 : hue_tab <= 6'd33;
			12'd2413 : hue_tab <= 6'd32;
			12'd2414 : hue_tab <= 6'd32;
			12'd2415 : hue_tab <= 6'd31;
			12'd2416 : hue_tab <= 6'd30;
			12'd2417 : hue_tab <= 6'd30;
			12'd2418 : hue_tab <= 6'd29;
			12'd2419 : hue_tab <= 6'd29;
			12'd2420 : hue_tab <= 6'd28;
			12'd2421 : hue_tab <= 6'd27;
			12'd2422 : hue_tab <= 6'd27;
			12'd2423 : hue_tab <= 6'd26;
			12'd2424 : hue_tab <= 6'd26;
			12'd2425 : hue_tab <= 6'd25;
			12'd2426 : hue_tab <= 6'd25;
			12'd2427 : hue_tab <= 6'd25;
			12'd2428 : hue_tab <= 6'd24;
			12'd2429 : hue_tab <= 6'd24;
			12'd2430 : hue_tab <= 6'd23;
			12'd2431 : hue_tab <= 6'd23;
			12'd2432 : hue_tab <= 6'd0;
			12'd2433 : hue_tab <= 6'd40;
			12'd2434 : hue_tab <= 6'd40;
			12'd2435 : hue_tab <= 6'd40;
			12'd2436 : hue_tab <= 6'd40;
			12'd2437 : hue_tab <= 6'd40;
			12'd2438 : hue_tab <= 6'd40;
			12'd2439 : hue_tab <= 6'd40;
			12'd2440 : hue_tab <= 6'd40;
			12'd2441 : hue_tab <= 6'd40;
			12'd2442 : hue_tab <= 6'd40;
			12'd2443 : hue_tab <= 6'd40;
			12'd2444 : hue_tab <= 6'd40;
			12'd2445 : hue_tab <= 6'd40;
			12'd2446 : hue_tab <= 6'd40;
			12'd2447 : hue_tab <= 6'd40;
			12'd2448 : hue_tab <= 6'd40;
			12'd2449 : hue_tab <= 6'd40;
			12'd2450 : hue_tab <= 6'd40;
			12'd2451 : hue_tab <= 6'd40;
			12'd2452 : hue_tab <= 6'd40;
			12'd2453 : hue_tab <= 6'd40;
			12'd2454 : hue_tab <= 6'd40;
			12'd2455 : hue_tab <= 6'd40;
			12'd2456 : hue_tab <= 6'd40;
			12'd2457 : hue_tab <= 6'd40;
			12'd2458 : hue_tab <= 6'd40;
			12'd2459 : hue_tab <= 6'd40;
			12'd2460 : hue_tab <= 6'd40;
			12'd2461 : hue_tab <= 6'd40;
			12'd2462 : hue_tab <= 6'd40;
			12'd2463 : hue_tab <= 6'd40;
			12'd2464 : hue_tab <= 6'd40;
			12'd2465 : hue_tab <= 6'd40;
			12'd2466 : hue_tab <= 6'd40;
			12'd2467 : hue_tab <= 6'd40;
			12'd2468 : hue_tab <= 6'd40;
			12'd2469 : hue_tab <= 6'd40;
			12'd2470 : hue_tab <= 6'd40;
			12'd2471 : hue_tab <= 6'd38;
			12'd2472 : hue_tab <= 6'd38;
			12'd2473 : hue_tab <= 6'd37;
			12'd2474 : hue_tab <= 6'd36;
			12'd2475 : hue_tab <= 6'd35;
			12'd2476 : hue_tab <= 6'd34;
			12'd2477 : hue_tab <= 6'd33;
			12'd2478 : hue_tab <= 6'd33;
			12'd2479 : hue_tab <= 6'd32;
			12'd2480 : hue_tab <= 6'd31;
			12'd2481 : hue_tab <= 6'd31;
			12'd2482 : hue_tab <= 6'd30;
			12'd2483 : hue_tab <= 6'd29;
			12'd2484 : hue_tab <= 6'd29;
			12'd2485 : hue_tab <= 6'd28;
			12'd2486 : hue_tab <= 6'd28;
			12'd2487 : hue_tab <= 6'd27;
			12'd2488 : hue_tab <= 6'd27;
			12'd2489 : hue_tab <= 6'd26;
			12'd2490 : hue_tab <= 6'd26;
			12'd2491 : hue_tab <= 6'd25;
			12'd2492 : hue_tab <= 6'd25;
			12'd2493 : hue_tab <= 6'd24;
			12'd2494 : hue_tab <= 6'd24;
			12'd2495 : hue_tab <= 6'd24;
			12'd2496 : hue_tab <= 6'd0;
			12'd2497 : hue_tab <= 6'd40;
			12'd2498 : hue_tab <= 6'd40;
			12'd2499 : hue_tab <= 6'd40;
			12'd2500 : hue_tab <= 6'd40;
			12'd2501 : hue_tab <= 6'd40;
			12'd2502 : hue_tab <= 6'd40;
			12'd2503 : hue_tab <= 6'd40;
			12'd2504 : hue_tab <= 6'd40;
			12'd2505 : hue_tab <= 6'd40;
			12'd2506 : hue_tab <= 6'd40;
			12'd2507 : hue_tab <= 6'd40;
			12'd2508 : hue_tab <= 6'd40;
			12'd2509 : hue_tab <= 6'd40;
			12'd2510 : hue_tab <= 6'd40;
			12'd2511 : hue_tab <= 6'd40;
			12'd2512 : hue_tab <= 6'd40;
			12'd2513 : hue_tab <= 6'd40;
			12'd2514 : hue_tab <= 6'd40;
			12'd2515 : hue_tab <= 6'd40;
			12'd2516 : hue_tab <= 6'd40;
			12'd2517 : hue_tab <= 6'd40;
			12'd2518 : hue_tab <= 6'd40;
			12'd2519 : hue_tab <= 6'd40;
			12'd2520 : hue_tab <= 6'd40;
			12'd2521 : hue_tab <= 6'd40;
			12'd2522 : hue_tab <= 6'd40;
			12'd2523 : hue_tab <= 6'd40;
			12'd2524 : hue_tab <= 6'd40;
			12'd2525 : hue_tab <= 6'd40;
			12'd2526 : hue_tab <= 6'd40;
			12'd2527 : hue_tab <= 6'd40;
			12'd2528 : hue_tab <= 6'd40;
			12'd2529 : hue_tab <= 6'd40;
			12'd2530 : hue_tab <= 6'd40;
			12'd2531 : hue_tab <= 6'd40;
			12'd2532 : hue_tab <= 6'd40;
			12'd2533 : hue_tab <= 6'd40;
			12'd2534 : hue_tab <= 6'd40;
			12'd2535 : hue_tab <= 6'd40;
			12'd2536 : hue_tab <= 6'd39;
			12'd2537 : hue_tab <= 6'd38;
			12'd2538 : hue_tab <= 6'd37;
			12'd2539 : hue_tab <= 6'd36;
			12'd2540 : hue_tab <= 6'd35;
			12'd2541 : hue_tab <= 6'd34;
			12'd2542 : hue_tab <= 6'd33;
			12'd2543 : hue_tab <= 6'd33;
			12'd2544 : hue_tab <= 6'd32;
			12'd2545 : hue_tab <= 6'd31;
			12'd2546 : hue_tab <= 6'd31;
			12'd2547 : hue_tab <= 6'd30;
			12'd2548 : hue_tab <= 6'd30;
			12'd2549 : hue_tab <= 6'd29;
			12'd2550 : hue_tab <= 6'd28;
			12'd2551 : hue_tab <= 6'd28;
			12'd2552 : hue_tab <= 6'd27;
			12'd2553 : hue_tab <= 6'd27;
			12'd2554 : hue_tab <= 6'd26;
			12'd2555 : hue_tab <= 6'd26;
			12'd2556 : hue_tab <= 6'd26;
			12'd2557 : hue_tab <= 6'd25;
			12'd2558 : hue_tab <= 6'd25;
			12'd2559 : hue_tab <= 6'd24;
			12'd2560 : hue_tab <= 6'd0;
			12'd2561 : hue_tab <= 6'd40;
			12'd2562 : hue_tab <= 6'd40;
			12'd2563 : hue_tab <= 6'd40;
			12'd2564 : hue_tab <= 6'd40;
			12'd2565 : hue_tab <= 6'd40;
			12'd2566 : hue_tab <= 6'd40;
			12'd2567 : hue_tab <= 6'd40;
			12'd2568 : hue_tab <= 6'd40;
			12'd2569 : hue_tab <= 6'd40;
			12'd2570 : hue_tab <= 6'd40;
			12'd2571 : hue_tab <= 6'd40;
			12'd2572 : hue_tab <= 6'd40;
			12'd2573 : hue_tab <= 6'd40;
			12'd2574 : hue_tab <= 6'd40;
			12'd2575 : hue_tab <= 6'd40;
			12'd2576 : hue_tab <= 6'd40;
			12'd2577 : hue_tab <= 6'd40;
			12'd2578 : hue_tab <= 6'd40;
			12'd2579 : hue_tab <= 6'd40;
			12'd2580 : hue_tab <= 6'd40;
			12'd2581 : hue_tab <= 6'd40;
			12'd2582 : hue_tab <= 6'd40;
			12'd2583 : hue_tab <= 6'd40;
			12'd2584 : hue_tab <= 6'd40;
			12'd2585 : hue_tab <= 6'd40;
			12'd2586 : hue_tab <= 6'd40;
			12'd2587 : hue_tab <= 6'd40;
			12'd2588 : hue_tab <= 6'd40;
			12'd2589 : hue_tab <= 6'd40;
			12'd2590 : hue_tab <= 6'd40;
			12'd2591 : hue_tab <= 6'd40;
			12'd2592 : hue_tab <= 6'd40;
			12'd2593 : hue_tab <= 6'd40;
			12'd2594 : hue_tab <= 6'd40;
			12'd2595 : hue_tab <= 6'd40;
			12'd2596 : hue_tab <= 6'd40;
			12'd2597 : hue_tab <= 6'd40;
			12'd2598 : hue_tab <= 6'd40;
			12'd2599 : hue_tab <= 6'd40;
			12'd2600 : hue_tab <= 6'd40;
			12'd2601 : hue_tab <= 6'd39;
			12'd2602 : hue_tab <= 6'd38;
			12'd2603 : hue_tab <= 6'd37;
			12'd2604 : hue_tab <= 6'd36;
			12'd2605 : hue_tab <= 6'd35;
			12'd2606 : hue_tab <= 6'd34;
			12'd2607 : hue_tab <= 6'd34;
			12'd2608 : hue_tab <= 6'd33;
			12'd2609 : hue_tab <= 6'd32;
			12'd2610 : hue_tab <= 6'd32;
			12'd2611 : hue_tab <= 6'd31;
			12'd2612 : hue_tab <= 6'd30;
			12'd2613 : hue_tab <= 6'd30;
			12'd2614 : hue_tab <= 6'd29;
			12'd2615 : hue_tab <= 6'd29;
			12'd2616 : hue_tab <= 6'd28;
			12'd2617 : hue_tab <= 6'd28;
			12'd2618 : hue_tab <= 6'd27;
			12'd2619 : hue_tab <= 6'd27;
			12'd2620 : hue_tab <= 6'd26;
			12'd2621 : hue_tab <= 6'd26;
			12'd2622 : hue_tab <= 6'd25;
			12'd2623 : hue_tab <= 6'd25;
			12'd2624 : hue_tab <= 6'd0;
			12'd2625 : hue_tab <= 6'd40;
			12'd2626 : hue_tab <= 6'd40;
			12'd2627 : hue_tab <= 6'd40;
			12'd2628 : hue_tab <= 6'd40;
			12'd2629 : hue_tab <= 6'd40;
			12'd2630 : hue_tab <= 6'd40;
			12'd2631 : hue_tab <= 6'd40;
			12'd2632 : hue_tab <= 6'd40;
			12'd2633 : hue_tab <= 6'd40;
			12'd2634 : hue_tab <= 6'd40;
			12'd2635 : hue_tab <= 6'd40;
			12'd2636 : hue_tab <= 6'd40;
			12'd2637 : hue_tab <= 6'd40;
			12'd2638 : hue_tab <= 6'd40;
			12'd2639 : hue_tab <= 6'd40;
			12'd2640 : hue_tab <= 6'd40;
			12'd2641 : hue_tab <= 6'd40;
			12'd2642 : hue_tab <= 6'd40;
			12'd2643 : hue_tab <= 6'd40;
			12'd2644 : hue_tab <= 6'd40;
			12'd2645 : hue_tab <= 6'd40;
			12'd2646 : hue_tab <= 6'd40;
			12'd2647 : hue_tab <= 6'd40;
			12'd2648 : hue_tab <= 6'd40;
			12'd2649 : hue_tab <= 6'd40;
			12'd2650 : hue_tab <= 6'd40;
			12'd2651 : hue_tab <= 6'd40;
			12'd2652 : hue_tab <= 6'd40;
			12'd2653 : hue_tab <= 6'd40;
			12'd2654 : hue_tab <= 6'd40;
			12'd2655 : hue_tab <= 6'd40;
			12'd2656 : hue_tab <= 6'd40;
			12'd2657 : hue_tab <= 6'd40;
			12'd2658 : hue_tab <= 6'd40;
			12'd2659 : hue_tab <= 6'd40;
			12'd2660 : hue_tab <= 6'd40;
			12'd2661 : hue_tab <= 6'd40;
			12'd2662 : hue_tab <= 6'd40;
			12'd2663 : hue_tab <= 6'd40;
			12'd2664 : hue_tab <= 6'd40;
			12'd2665 : hue_tab <= 6'd40;
			12'd2666 : hue_tab <= 6'd39;
			12'd2667 : hue_tab <= 6'd38;
			12'd2668 : hue_tab <= 6'd37;
			12'd2669 : hue_tab <= 6'd36;
			12'd2670 : hue_tab <= 6'd35;
			12'd2671 : hue_tab <= 6'd34;
			12'd2672 : hue_tab <= 6'd34;
			12'd2673 : hue_tab <= 6'd33;
			12'd2674 : hue_tab <= 6'd32;
			12'd2675 : hue_tab <= 6'd32;
			12'd2676 : hue_tab <= 6'd31;
			12'd2677 : hue_tab <= 6'd30;
			12'd2678 : hue_tab <= 6'd30;
			12'd2679 : hue_tab <= 6'd29;
			12'd2680 : hue_tab <= 6'd29;
			12'd2681 : hue_tab <= 6'd28;
			12'd2682 : hue_tab <= 6'd28;
			12'd2683 : hue_tab <= 6'd27;
			12'd2684 : hue_tab <= 6'd27;
			12'd2685 : hue_tab <= 6'd26;
			12'd2686 : hue_tab <= 6'd26;
			12'd2687 : hue_tab <= 6'd26;
			12'd2688 : hue_tab <= 6'd0;
			12'd2689 : hue_tab <= 6'd40;
			12'd2690 : hue_tab <= 6'd40;
			12'd2691 : hue_tab <= 6'd40;
			12'd2692 : hue_tab <= 6'd40;
			12'd2693 : hue_tab <= 6'd40;
			12'd2694 : hue_tab <= 6'd40;
			12'd2695 : hue_tab <= 6'd40;
			12'd2696 : hue_tab <= 6'd40;
			12'd2697 : hue_tab <= 6'd40;
			12'd2698 : hue_tab <= 6'd40;
			12'd2699 : hue_tab <= 6'd40;
			12'd2700 : hue_tab <= 6'd40;
			12'd2701 : hue_tab <= 6'd40;
			12'd2702 : hue_tab <= 6'd40;
			12'd2703 : hue_tab <= 6'd40;
			12'd2704 : hue_tab <= 6'd40;
			12'd2705 : hue_tab <= 6'd40;
			12'd2706 : hue_tab <= 6'd40;
			12'd2707 : hue_tab <= 6'd40;
			12'd2708 : hue_tab <= 6'd40;
			12'd2709 : hue_tab <= 6'd40;
			12'd2710 : hue_tab <= 6'd40;
			12'd2711 : hue_tab <= 6'd40;
			12'd2712 : hue_tab <= 6'd40;
			12'd2713 : hue_tab <= 6'd40;
			12'd2714 : hue_tab <= 6'd40;
			12'd2715 : hue_tab <= 6'd40;
			12'd2716 : hue_tab <= 6'd40;
			12'd2717 : hue_tab <= 6'd40;
			12'd2718 : hue_tab <= 6'd40;
			12'd2719 : hue_tab <= 6'd40;
			12'd2720 : hue_tab <= 6'd40;
			12'd2721 : hue_tab <= 6'd40;
			12'd2722 : hue_tab <= 6'd40;
			12'd2723 : hue_tab <= 6'd40;
			12'd2724 : hue_tab <= 6'd40;
			12'd2725 : hue_tab <= 6'd40;
			12'd2726 : hue_tab <= 6'd40;
			12'd2727 : hue_tab <= 6'd40;
			12'd2728 : hue_tab <= 6'd40;
			12'd2729 : hue_tab <= 6'd40;
			12'd2730 : hue_tab <= 6'd40;
			12'd2731 : hue_tab <= 6'd39;
			12'd2732 : hue_tab <= 6'd38;
			12'd2733 : hue_tab <= 6'd37;
			12'd2734 : hue_tab <= 6'd36;
			12'd2735 : hue_tab <= 6'd35;
			12'd2736 : hue_tab <= 6'd35;
			12'd2737 : hue_tab <= 6'd34;
			12'd2738 : hue_tab <= 6'd33;
			12'd2739 : hue_tab <= 6'd32;
			12'd2740 : hue_tab <= 6'd32;
			12'd2741 : hue_tab <= 6'd31;
			12'd2742 : hue_tab <= 6'd31;
			12'd2743 : hue_tab <= 6'd30;
			12'd2744 : hue_tab <= 6'd30;
			12'd2745 : hue_tab <= 6'd29;
			12'd2746 : hue_tab <= 6'd28;
			12'd2747 : hue_tab <= 6'd28;
			12'd2748 : hue_tab <= 6'd28;
			12'd2749 : hue_tab <= 6'd27;
			12'd2750 : hue_tab <= 6'd27;
			12'd2751 : hue_tab <= 6'd26;
			12'd2752 : hue_tab <= 6'd0;
			12'd2753 : hue_tab <= 6'd40;
			12'd2754 : hue_tab <= 6'd40;
			12'd2755 : hue_tab <= 6'd40;
			12'd2756 : hue_tab <= 6'd40;
			12'd2757 : hue_tab <= 6'd40;
			12'd2758 : hue_tab <= 6'd40;
			12'd2759 : hue_tab <= 6'd40;
			12'd2760 : hue_tab <= 6'd40;
			12'd2761 : hue_tab <= 6'd40;
			12'd2762 : hue_tab <= 6'd40;
			12'd2763 : hue_tab <= 6'd40;
			12'd2764 : hue_tab <= 6'd40;
			12'd2765 : hue_tab <= 6'd40;
			12'd2766 : hue_tab <= 6'd40;
			12'd2767 : hue_tab <= 6'd40;
			12'd2768 : hue_tab <= 6'd40;
			12'd2769 : hue_tab <= 6'd40;
			12'd2770 : hue_tab <= 6'd40;
			12'd2771 : hue_tab <= 6'd40;
			12'd2772 : hue_tab <= 6'd40;
			12'd2773 : hue_tab <= 6'd40;
			12'd2774 : hue_tab <= 6'd40;
			12'd2775 : hue_tab <= 6'd40;
			12'd2776 : hue_tab <= 6'd40;
			12'd2777 : hue_tab <= 6'd40;
			12'd2778 : hue_tab <= 6'd40;
			12'd2779 : hue_tab <= 6'd40;
			12'd2780 : hue_tab <= 6'd40;
			12'd2781 : hue_tab <= 6'd40;
			12'd2782 : hue_tab <= 6'd40;
			12'd2783 : hue_tab <= 6'd40;
			12'd2784 : hue_tab <= 6'd40;
			12'd2785 : hue_tab <= 6'd40;
			12'd2786 : hue_tab <= 6'd40;
			12'd2787 : hue_tab <= 6'd40;
			12'd2788 : hue_tab <= 6'd40;
			12'd2789 : hue_tab <= 6'd40;
			12'd2790 : hue_tab <= 6'd40;
			12'd2791 : hue_tab <= 6'd40;
			12'd2792 : hue_tab <= 6'd40;
			12'd2793 : hue_tab <= 6'd40;
			12'd2794 : hue_tab <= 6'd40;
			12'd2795 : hue_tab <= 6'd40;
			12'd2796 : hue_tab <= 6'd39;
			12'd2797 : hue_tab <= 6'd38;
			12'd2798 : hue_tab <= 6'd37;
			12'd2799 : hue_tab <= 6'd36;
			12'd2800 : hue_tab <= 6'd35;
			12'd2801 : hue_tab <= 6'd35;
			12'd2802 : hue_tab <= 6'd34;
			12'd2803 : hue_tab <= 6'd33;
			12'd2804 : hue_tab <= 6'd33;
			12'd2805 : hue_tab <= 6'd32;
			12'd2806 : hue_tab <= 6'd31;
			12'd2807 : hue_tab <= 6'd31;
			12'd2808 : hue_tab <= 6'd30;
			12'd2809 : hue_tab <= 6'd30;
			12'd2810 : hue_tab <= 6'd29;
			12'd2811 : hue_tab <= 6'd29;
			12'd2812 : hue_tab <= 6'd28;
			12'd2813 : hue_tab <= 6'd28;
			12'd2814 : hue_tab <= 6'd27;
			12'd2815 : hue_tab <= 6'd27;
			12'd2816 : hue_tab <= 6'd0;
			12'd2817 : hue_tab <= 6'd40;
			12'd2818 : hue_tab <= 6'd40;
			12'd2819 : hue_tab <= 6'd40;
			12'd2820 : hue_tab <= 6'd40;
			12'd2821 : hue_tab <= 6'd40;
			12'd2822 : hue_tab <= 6'd40;
			12'd2823 : hue_tab <= 6'd40;
			12'd2824 : hue_tab <= 6'd40;
			12'd2825 : hue_tab <= 6'd40;
			12'd2826 : hue_tab <= 6'd40;
			12'd2827 : hue_tab <= 6'd40;
			12'd2828 : hue_tab <= 6'd40;
			12'd2829 : hue_tab <= 6'd40;
			12'd2830 : hue_tab <= 6'd40;
			12'd2831 : hue_tab <= 6'd40;
			12'd2832 : hue_tab <= 6'd40;
			12'd2833 : hue_tab <= 6'd40;
			12'd2834 : hue_tab <= 6'd40;
			12'd2835 : hue_tab <= 6'd40;
			12'd2836 : hue_tab <= 6'd40;
			12'd2837 : hue_tab <= 6'd40;
			12'd2838 : hue_tab <= 6'd40;
			12'd2839 : hue_tab <= 6'd40;
			12'd2840 : hue_tab <= 6'd40;
			12'd2841 : hue_tab <= 6'd40;
			12'd2842 : hue_tab <= 6'd40;
			12'd2843 : hue_tab <= 6'd40;
			12'd2844 : hue_tab <= 6'd40;
			12'd2845 : hue_tab <= 6'd40;
			12'd2846 : hue_tab <= 6'd40;
			12'd2847 : hue_tab <= 6'd40;
			12'd2848 : hue_tab <= 6'd40;
			12'd2849 : hue_tab <= 6'd40;
			12'd2850 : hue_tab <= 6'd40;
			12'd2851 : hue_tab <= 6'd40;
			12'd2852 : hue_tab <= 6'd40;
			12'd2853 : hue_tab <= 6'd40;
			12'd2854 : hue_tab <= 6'd40;
			12'd2855 : hue_tab <= 6'd40;
			12'd2856 : hue_tab <= 6'd40;
			12'd2857 : hue_tab <= 6'd40;
			12'd2858 : hue_tab <= 6'd40;
			12'd2859 : hue_tab <= 6'd40;
			12'd2860 : hue_tab <= 6'd40;
			12'd2861 : hue_tab <= 6'd39;
			12'd2862 : hue_tab <= 6'd38;
			12'd2863 : hue_tab <= 6'd37;
			12'd2864 : hue_tab <= 6'd36;
			12'd2865 : hue_tab <= 6'd35;
			12'd2866 : hue_tab <= 6'd35;
			12'd2867 : hue_tab <= 6'd34;
			12'd2868 : hue_tab <= 6'd33;
			12'd2869 : hue_tab <= 6'd33;
			12'd2870 : hue_tab <= 6'd32;
			12'd2871 : hue_tab <= 6'd32;
			12'd2872 : hue_tab <= 6'd31;
			12'd2873 : hue_tab <= 6'd30;
			12'd2874 : hue_tab <= 6'd30;
			12'd2875 : hue_tab <= 6'd29;
			12'd2876 : hue_tab <= 6'd29;
			12'd2877 : hue_tab <= 6'd28;
			12'd2878 : hue_tab <= 6'd28;
			12'd2879 : hue_tab <= 6'd27;
			12'd2880 : hue_tab <= 6'd0;
			12'd2881 : hue_tab <= 6'd40;
			12'd2882 : hue_tab <= 6'd40;
			12'd2883 : hue_tab <= 6'd40;
			12'd2884 : hue_tab <= 6'd40;
			12'd2885 : hue_tab <= 6'd40;
			12'd2886 : hue_tab <= 6'd40;
			12'd2887 : hue_tab <= 6'd40;
			12'd2888 : hue_tab <= 6'd40;
			12'd2889 : hue_tab <= 6'd40;
			12'd2890 : hue_tab <= 6'd40;
			12'd2891 : hue_tab <= 6'd40;
			12'd2892 : hue_tab <= 6'd40;
			12'd2893 : hue_tab <= 6'd40;
			12'd2894 : hue_tab <= 6'd40;
			12'd2895 : hue_tab <= 6'd40;
			12'd2896 : hue_tab <= 6'd40;
			12'd2897 : hue_tab <= 6'd40;
			12'd2898 : hue_tab <= 6'd40;
			12'd2899 : hue_tab <= 6'd40;
			12'd2900 : hue_tab <= 6'd40;
			12'd2901 : hue_tab <= 6'd40;
			12'd2902 : hue_tab <= 6'd40;
			12'd2903 : hue_tab <= 6'd40;
			12'd2904 : hue_tab <= 6'd40;
			12'd2905 : hue_tab <= 6'd40;
			12'd2906 : hue_tab <= 6'd40;
			12'd2907 : hue_tab <= 6'd40;
			12'd2908 : hue_tab <= 6'd40;
			12'd2909 : hue_tab <= 6'd40;
			12'd2910 : hue_tab <= 6'd40;
			12'd2911 : hue_tab <= 6'd40;
			12'd2912 : hue_tab <= 6'd40;
			12'd2913 : hue_tab <= 6'd40;
			12'd2914 : hue_tab <= 6'd40;
			12'd2915 : hue_tab <= 6'd40;
			12'd2916 : hue_tab <= 6'd40;
			12'd2917 : hue_tab <= 6'd40;
			12'd2918 : hue_tab <= 6'd40;
			12'd2919 : hue_tab <= 6'd40;
			12'd2920 : hue_tab <= 6'd40;
			12'd2921 : hue_tab <= 6'd40;
			12'd2922 : hue_tab <= 6'd40;
			12'd2923 : hue_tab <= 6'd40;
			12'd2924 : hue_tab <= 6'd40;
			12'd2925 : hue_tab <= 6'd40;
			12'd2926 : hue_tab <= 6'd39;
			12'd2927 : hue_tab <= 6'd38;
			12'd2928 : hue_tab <= 6'd37;
			12'd2929 : hue_tab <= 6'd36;
			12'd2930 : hue_tab <= 6'd36;
			12'd2931 : hue_tab <= 6'd35;
			12'd2932 : hue_tab <= 6'd34;
			12'd2933 : hue_tab <= 6'd33;
			12'd2934 : hue_tab <= 6'd33;
			12'd2935 : hue_tab <= 6'd32;
			12'd2936 : hue_tab <= 6'd32;
			12'd2937 : hue_tab <= 6'd31;
			12'd2938 : hue_tab <= 6'd31;
			12'd2939 : hue_tab <= 6'd30;
			12'd2940 : hue_tab <= 6'd30;
			12'd2941 : hue_tab <= 6'd29;
			12'd2942 : hue_tab <= 6'd29;
			12'd2943 : hue_tab <= 6'd28;
			12'd2944 : hue_tab <= 6'd0;
			12'd2945 : hue_tab <= 6'd40;
			12'd2946 : hue_tab <= 6'd40;
			12'd2947 : hue_tab <= 6'd40;
			12'd2948 : hue_tab <= 6'd40;
			12'd2949 : hue_tab <= 6'd40;
			12'd2950 : hue_tab <= 6'd40;
			12'd2951 : hue_tab <= 6'd40;
			12'd2952 : hue_tab <= 6'd40;
			12'd2953 : hue_tab <= 6'd40;
			12'd2954 : hue_tab <= 6'd40;
			12'd2955 : hue_tab <= 6'd40;
			12'd2956 : hue_tab <= 6'd40;
			12'd2957 : hue_tab <= 6'd40;
			12'd2958 : hue_tab <= 6'd40;
			12'd2959 : hue_tab <= 6'd40;
			12'd2960 : hue_tab <= 6'd40;
			12'd2961 : hue_tab <= 6'd40;
			12'd2962 : hue_tab <= 6'd40;
			12'd2963 : hue_tab <= 6'd40;
			12'd2964 : hue_tab <= 6'd40;
			12'd2965 : hue_tab <= 6'd40;
			12'd2966 : hue_tab <= 6'd40;
			12'd2967 : hue_tab <= 6'd40;
			12'd2968 : hue_tab <= 6'd40;
			12'd2969 : hue_tab <= 6'd40;
			12'd2970 : hue_tab <= 6'd40;
			12'd2971 : hue_tab <= 6'd40;
			12'd2972 : hue_tab <= 6'd40;
			12'd2973 : hue_tab <= 6'd40;
			12'd2974 : hue_tab <= 6'd40;
			12'd2975 : hue_tab <= 6'd40;
			12'd2976 : hue_tab <= 6'd40;
			12'd2977 : hue_tab <= 6'd40;
			12'd2978 : hue_tab <= 6'd40;
			12'd2979 : hue_tab <= 6'd40;
			12'd2980 : hue_tab <= 6'd40;
			12'd2981 : hue_tab <= 6'd40;
			12'd2982 : hue_tab <= 6'd40;
			12'd2983 : hue_tab <= 6'd40;
			12'd2984 : hue_tab <= 6'd40;
			12'd2985 : hue_tab <= 6'd40;
			12'd2986 : hue_tab <= 6'd40;
			12'd2987 : hue_tab <= 6'd40;
			12'd2988 : hue_tab <= 6'd40;
			12'd2989 : hue_tab <= 6'd40;
			12'd2990 : hue_tab <= 6'd40;
			12'd2991 : hue_tab <= 6'd39;
			12'd2992 : hue_tab <= 6'd38;
			12'd2993 : hue_tab <= 6'd37;
			12'd2994 : hue_tab <= 6'd36;
			12'd2995 : hue_tab <= 6'd36;
			12'd2996 : hue_tab <= 6'd35;
			12'd2997 : hue_tab <= 6'd34;
			12'd2998 : hue_tab <= 6'd34;
			12'd2999 : hue_tab <= 6'd33;
			12'd3000 : hue_tab <= 6'd32;
			12'd3001 : hue_tab <= 6'd32;
			12'd3002 : hue_tab <= 6'd31;
			12'd3003 : hue_tab <= 6'd31;
			12'd3004 : hue_tab <= 6'd30;
			12'd3005 : hue_tab <= 6'd30;
			12'd3006 : hue_tab <= 6'd29;
			12'd3007 : hue_tab <= 6'd29;
			12'd3008 : hue_tab <= 6'd0;
			12'd3009 : hue_tab <= 6'd40;
			12'd3010 : hue_tab <= 6'd40;
			12'd3011 : hue_tab <= 6'd40;
			12'd3012 : hue_tab <= 6'd40;
			12'd3013 : hue_tab <= 6'd40;
			12'd3014 : hue_tab <= 6'd40;
			12'd3015 : hue_tab <= 6'd40;
			12'd3016 : hue_tab <= 6'd40;
			12'd3017 : hue_tab <= 6'd40;
			12'd3018 : hue_tab <= 6'd40;
			12'd3019 : hue_tab <= 6'd40;
			12'd3020 : hue_tab <= 6'd40;
			12'd3021 : hue_tab <= 6'd40;
			12'd3022 : hue_tab <= 6'd40;
			12'd3023 : hue_tab <= 6'd40;
			12'd3024 : hue_tab <= 6'd40;
			12'd3025 : hue_tab <= 6'd40;
			12'd3026 : hue_tab <= 6'd40;
			12'd3027 : hue_tab <= 6'd40;
			12'd3028 : hue_tab <= 6'd40;
			12'd3029 : hue_tab <= 6'd40;
			12'd3030 : hue_tab <= 6'd40;
			12'd3031 : hue_tab <= 6'd40;
			12'd3032 : hue_tab <= 6'd40;
			12'd3033 : hue_tab <= 6'd40;
			12'd3034 : hue_tab <= 6'd40;
			12'd3035 : hue_tab <= 6'd40;
			12'd3036 : hue_tab <= 6'd40;
			12'd3037 : hue_tab <= 6'd40;
			12'd3038 : hue_tab <= 6'd40;
			12'd3039 : hue_tab <= 6'd40;
			12'd3040 : hue_tab <= 6'd40;
			12'd3041 : hue_tab <= 6'd40;
			12'd3042 : hue_tab <= 6'd40;
			12'd3043 : hue_tab <= 6'd40;
			12'd3044 : hue_tab <= 6'd40;
			12'd3045 : hue_tab <= 6'd40;
			12'd3046 : hue_tab <= 6'd40;
			12'd3047 : hue_tab <= 6'd40;
			12'd3048 : hue_tab <= 6'd40;
			12'd3049 : hue_tab <= 6'd40;
			12'd3050 : hue_tab <= 6'd40;
			12'd3051 : hue_tab <= 6'd40;
			12'd3052 : hue_tab <= 6'd40;
			12'd3053 : hue_tab <= 6'd40;
			12'd3054 : hue_tab <= 6'd40;
			12'd3055 : hue_tab <= 6'd40;
			12'd3056 : hue_tab <= 6'd39;
			12'd3057 : hue_tab <= 6'd38;
			12'd3058 : hue_tab <= 6'd37;
			12'd3059 : hue_tab <= 6'd36;
			12'd3060 : hue_tab <= 6'd36;
			12'd3061 : hue_tab <= 6'd35;
			12'd3062 : hue_tab <= 6'd34;
			12'd3063 : hue_tab <= 6'd34;
			12'd3064 : hue_tab <= 6'd33;
			12'd3065 : hue_tab <= 6'd32;
			12'd3066 : hue_tab <= 6'd32;
			12'd3067 : hue_tab <= 6'd31;
			12'd3068 : hue_tab <= 6'd31;
			12'd3069 : hue_tab <= 6'd30;
			12'd3070 : hue_tab <= 6'd30;
			12'd3071 : hue_tab <= 6'd29;
			12'd3072 : hue_tab <= 6'd0;
			12'd3073 : hue_tab <= 6'd40;
			12'd3074 : hue_tab <= 6'd40;
			12'd3075 : hue_tab <= 6'd40;
			12'd3076 : hue_tab <= 6'd40;
			12'd3077 : hue_tab <= 6'd40;
			12'd3078 : hue_tab <= 6'd40;
			12'd3079 : hue_tab <= 6'd40;
			12'd3080 : hue_tab <= 6'd40;
			12'd3081 : hue_tab <= 6'd40;
			12'd3082 : hue_tab <= 6'd40;
			12'd3083 : hue_tab <= 6'd40;
			12'd3084 : hue_tab <= 6'd40;
			12'd3085 : hue_tab <= 6'd40;
			12'd3086 : hue_tab <= 6'd40;
			12'd3087 : hue_tab <= 6'd40;
			12'd3088 : hue_tab <= 6'd40;
			12'd3089 : hue_tab <= 6'd40;
			12'd3090 : hue_tab <= 6'd40;
			12'd3091 : hue_tab <= 6'd40;
			12'd3092 : hue_tab <= 6'd40;
			12'd3093 : hue_tab <= 6'd40;
			12'd3094 : hue_tab <= 6'd40;
			12'd3095 : hue_tab <= 6'd40;
			12'd3096 : hue_tab <= 6'd40;
			12'd3097 : hue_tab <= 6'd40;
			12'd3098 : hue_tab <= 6'd40;
			12'd3099 : hue_tab <= 6'd40;
			12'd3100 : hue_tab <= 6'd40;
			12'd3101 : hue_tab <= 6'd40;
			12'd3102 : hue_tab <= 6'd40;
			12'd3103 : hue_tab <= 6'd40;
			12'd3104 : hue_tab <= 6'd40;
			12'd3105 : hue_tab <= 6'd40;
			12'd3106 : hue_tab <= 6'd40;
			12'd3107 : hue_tab <= 6'd40;
			12'd3108 : hue_tab <= 6'd40;
			12'd3109 : hue_tab <= 6'd40;
			12'd3110 : hue_tab <= 6'd40;
			12'd3111 : hue_tab <= 6'd40;
			12'd3112 : hue_tab <= 6'd40;
			12'd3113 : hue_tab <= 6'd40;
			12'd3114 : hue_tab <= 6'd40;
			12'd3115 : hue_tab <= 6'd40;
			12'd3116 : hue_tab <= 6'd40;
			12'd3117 : hue_tab <= 6'd40;
			12'd3118 : hue_tab <= 6'd40;
			12'd3119 : hue_tab <= 6'd40;
			12'd3120 : hue_tab <= 6'd40;
			12'd3121 : hue_tab <= 6'd39;
			12'd3122 : hue_tab <= 6'd38;
			12'd3123 : hue_tab <= 6'd37;
			12'd3124 : hue_tab <= 6'd36;
			12'd3125 : hue_tab <= 6'd36;
			12'd3126 : hue_tab <= 6'd35;
			12'd3127 : hue_tab <= 6'd34;
			12'd3128 : hue_tab <= 6'd34;
			12'd3129 : hue_tab <= 6'd33;
			12'd3130 : hue_tab <= 6'd33;
			12'd3131 : hue_tab <= 6'd32;
			12'd3132 : hue_tab <= 6'd32;
			12'd3133 : hue_tab <= 6'd31;
			12'd3134 : hue_tab <= 6'd30;
			12'd3135 : hue_tab <= 6'd30;
			12'd3136 : hue_tab <= 6'd0;
			12'd3137 : hue_tab <= 6'd40;
			12'd3138 : hue_tab <= 6'd40;
			12'd3139 : hue_tab <= 6'd40;
			12'd3140 : hue_tab <= 6'd40;
			12'd3141 : hue_tab <= 6'd40;
			12'd3142 : hue_tab <= 6'd40;
			12'd3143 : hue_tab <= 6'd40;
			12'd3144 : hue_tab <= 6'd40;
			12'd3145 : hue_tab <= 6'd40;
			12'd3146 : hue_tab <= 6'd40;
			12'd3147 : hue_tab <= 6'd40;
			12'd3148 : hue_tab <= 6'd40;
			12'd3149 : hue_tab <= 6'd40;
			12'd3150 : hue_tab <= 6'd40;
			12'd3151 : hue_tab <= 6'd40;
			12'd3152 : hue_tab <= 6'd40;
			12'd3153 : hue_tab <= 6'd40;
			12'd3154 : hue_tab <= 6'd40;
			12'd3155 : hue_tab <= 6'd40;
			12'd3156 : hue_tab <= 6'd40;
			12'd3157 : hue_tab <= 6'd40;
			12'd3158 : hue_tab <= 6'd40;
			12'd3159 : hue_tab <= 6'd40;
			12'd3160 : hue_tab <= 6'd40;
			12'd3161 : hue_tab <= 6'd40;
			12'd3162 : hue_tab <= 6'd40;
			12'd3163 : hue_tab <= 6'd40;
			12'd3164 : hue_tab <= 6'd40;
			12'd3165 : hue_tab <= 6'd40;
			12'd3166 : hue_tab <= 6'd40;
			12'd3167 : hue_tab <= 6'd40;
			12'd3168 : hue_tab <= 6'd40;
			12'd3169 : hue_tab <= 6'd40;
			12'd3170 : hue_tab <= 6'd40;
			12'd3171 : hue_tab <= 6'd40;
			12'd3172 : hue_tab <= 6'd40;
			12'd3173 : hue_tab <= 6'd40;
			12'd3174 : hue_tab <= 6'd40;
			12'd3175 : hue_tab <= 6'd40;
			12'd3176 : hue_tab <= 6'd40;
			12'd3177 : hue_tab <= 6'd40;
			12'd3178 : hue_tab <= 6'd40;
			12'd3179 : hue_tab <= 6'd40;
			12'd3180 : hue_tab <= 6'd40;
			12'd3181 : hue_tab <= 6'd40;
			12'd3182 : hue_tab <= 6'd40;
			12'd3183 : hue_tab <= 6'd40;
			12'd3184 : hue_tab <= 6'd40;
			12'd3185 : hue_tab <= 6'd40;
			12'd3186 : hue_tab <= 6'd39;
			12'd3187 : hue_tab <= 6'd38;
			12'd3188 : hue_tab <= 6'd37;
			12'd3189 : hue_tab <= 6'd36;
			12'd3190 : hue_tab <= 6'd36;
			12'd3191 : hue_tab <= 6'd35;
			12'd3192 : hue_tab <= 6'd35;
			12'd3193 : hue_tab <= 6'd34;
			12'd3194 : hue_tab <= 6'd33;
			12'd3195 : hue_tab <= 6'd33;
			12'd3196 : hue_tab <= 6'd32;
			12'd3197 : hue_tab <= 6'd32;
			12'd3198 : hue_tab <= 6'd31;
			12'd3199 : hue_tab <= 6'd31;
			12'd3200 : hue_tab <= 6'd0;
			12'd3201 : hue_tab <= 6'd40;
			12'd3202 : hue_tab <= 6'd40;
			12'd3203 : hue_tab <= 6'd40;
			12'd3204 : hue_tab <= 6'd40;
			12'd3205 : hue_tab <= 6'd40;
			12'd3206 : hue_tab <= 6'd40;
			12'd3207 : hue_tab <= 6'd40;
			12'd3208 : hue_tab <= 6'd40;
			12'd3209 : hue_tab <= 6'd40;
			12'd3210 : hue_tab <= 6'd40;
			12'd3211 : hue_tab <= 6'd40;
			12'd3212 : hue_tab <= 6'd40;
			12'd3213 : hue_tab <= 6'd40;
			12'd3214 : hue_tab <= 6'd40;
			12'd3215 : hue_tab <= 6'd40;
			12'd3216 : hue_tab <= 6'd40;
			12'd3217 : hue_tab <= 6'd40;
			12'd3218 : hue_tab <= 6'd40;
			12'd3219 : hue_tab <= 6'd40;
			12'd3220 : hue_tab <= 6'd40;
			12'd3221 : hue_tab <= 6'd40;
			12'd3222 : hue_tab <= 6'd40;
			12'd3223 : hue_tab <= 6'd40;
			12'd3224 : hue_tab <= 6'd40;
			12'd3225 : hue_tab <= 6'd40;
			12'd3226 : hue_tab <= 6'd40;
			12'd3227 : hue_tab <= 6'd40;
			12'd3228 : hue_tab <= 6'd40;
			12'd3229 : hue_tab <= 6'd40;
			12'd3230 : hue_tab <= 6'd40;
			12'd3231 : hue_tab <= 6'd40;
			12'd3232 : hue_tab <= 6'd40;
			12'd3233 : hue_tab <= 6'd40;
			12'd3234 : hue_tab <= 6'd40;
			12'd3235 : hue_tab <= 6'd40;
			12'd3236 : hue_tab <= 6'd40;
			12'd3237 : hue_tab <= 6'd40;
			12'd3238 : hue_tab <= 6'd40;
			12'd3239 : hue_tab <= 6'd40;
			12'd3240 : hue_tab <= 6'd40;
			12'd3241 : hue_tab <= 6'd40;
			12'd3242 : hue_tab <= 6'd40;
			12'd3243 : hue_tab <= 6'd40;
			12'd3244 : hue_tab <= 6'd40;
			12'd3245 : hue_tab <= 6'd40;
			12'd3246 : hue_tab <= 6'd40;
			12'd3247 : hue_tab <= 6'd40;
			12'd3248 : hue_tab <= 6'd40;
			12'd3249 : hue_tab <= 6'd40;
			12'd3250 : hue_tab <= 6'd40;
			12'd3251 : hue_tab <= 6'd39;
			12'd3252 : hue_tab <= 6'd38;
			12'd3253 : hue_tab <= 6'd37;
			12'd3254 : hue_tab <= 6'd37;
			12'd3255 : hue_tab <= 6'd36;
			12'd3256 : hue_tab <= 6'd35;
			12'd3257 : hue_tab <= 6'd35;
			12'd3258 : hue_tab <= 6'd34;
			12'd3259 : hue_tab <= 6'd33;
			12'd3260 : hue_tab <= 6'd33;
			12'd3261 : hue_tab <= 6'd32;
			12'd3262 : hue_tab <= 6'd32;
			12'd3263 : hue_tab <= 6'd31;
			12'd3264 : hue_tab <= 6'd0;
			12'd3265 : hue_tab <= 6'd40;
			12'd3266 : hue_tab <= 6'd40;
			12'd3267 : hue_tab <= 6'd40;
			12'd3268 : hue_tab <= 6'd40;
			12'd3269 : hue_tab <= 6'd40;
			12'd3270 : hue_tab <= 6'd40;
			12'd3271 : hue_tab <= 6'd40;
			12'd3272 : hue_tab <= 6'd40;
			12'd3273 : hue_tab <= 6'd40;
			12'd3274 : hue_tab <= 6'd40;
			12'd3275 : hue_tab <= 6'd40;
			12'd3276 : hue_tab <= 6'd40;
			12'd3277 : hue_tab <= 6'd40;
			12'd3278 : hue_tab <= 6'd40;
			12'd3279 : hue_tab <= 6'd40;
			12'd3280 : hue_tab <= 6'd40;
			12'd3281 : hue_tab <= 6'd40;
			12'd3282 : hue_tab <= 6'd40;
			12'd3283 : hue_tab <= 6'd40;
			12'd3284 : hue_tab <= 6'd40;
			12'd3285 : hue_tab <= 6'd40;
			12'd3286 : hue_tab <= 6'd40;
			12'd3287 : hue_tab <= 6'd40;
			12'd3288 : hue_tab <= 6'd40;
			12'd3289 : hue_tab <= 6'd40;
			12'd3290 : hue_tab <= 6'd40;
			12'd3291 : hue_tab <= 6'd40;
			12'd3292 : hue_tab <= 6'd40;
			12'd3293 : hue_tab <= 6'd40;
			12'd3294 : hue_tab <= 6'd40;
			12'd3295 : hue_tab <= 6'd40;
			12'd3296 : hue_tab <= 6'd40;
			12'd3297 : hue_tab <= 6'd40;
			12'd3298 : hue_tab <= 6'd40;
			12'd3299 : hue_tab <= 6'd40;
			12'd3300 : hue_tab <= 6'd40;
			12'd3301 : hue_tab <= 6'd40;
			12'd3302 : hue_tab <= 6'd40;
			12'd3303 : hue_tab <= 6'd40;
			12'd3304 : hue_tab <= 6'd40;
			12'd3305 : hue_tab <= 6'd40;
			12'd3306 : hue_tab <= 6'd40;
			12'd3307 : hue_tab <= 6'd40;
			12'd3308 : hue_tab <= 6'd40;
			12'd3309 : hue_tab <= 6'd40;
			12'd3310 : hue_tab <= 6'd40;
			12'd3311 : hue_tab <= 6'd40;
			12'd3312 : hue_tab <= 6'd40;
			12'd3313 : hue_tab <= 6'd40;
			12'd3314 : hue_tab <= 6'd40;
			12'd3315 : hue_tab <= 6'd40;
			12'd3316 : hue_tab <= 6'd39;
			12'd3317 : hue_tab <= 6'd38;
			12'd3318 : hue_tab <= 6'd37;
			12'd3319 : hue_tab <= 6'd37;
			12'd3320 : hue_tab <= 6'd36;
			12'd3321 : hue_tab <= 6'd35;
			12'd3322 : hue_tab <= 6'd35;
			12'd3323 : hue_tab <= 6'd34;
			12'd3324 : hue_tab <= 6'd34;
			12'd3325 : hue_tab <= 6'd33;
			12'd3326 : hue_tab <= 6'd32;
			12'd3327 : hue_tab <= 6'd32;
			12'd3328 : hue_tab <= 6'd0;
			12'd3329 : hue_tab <= 6'd40;
			12'd3330 : hue_tab <= 6'd40;
			12'd3331 : hue_tab <= 6'd40;
			12'd3332 : hue_tab <= 6'd40;
			12'd3333 : hue_tab <= 6'd40;
			12'd3334 : hue_tab <= 6'd40;
			12'd3335 : hue_tab <= 6'd40;
			12'd3336 : hue_tab <= 6'd40;
			12'd3337 : hue_tab <= 6'd40;
			12'd3338 : hue_tab <= 6'd40;
			12'd3339 : hue_tab <= 6'd40;
			12'd3340 : hue_tab <= 6'd40;
			12'd3341 : hue_tab <= 6'd40;
			12'd3342 : hue_tab <= 6'd40;
			12'd3343 : hue_tab <= 6'd40;
			12'd3344 : hue_tab <= 6'd40;
			12'd3345 : hue_tab <= 6'd40;
			12'd3346 : hue_tab <= 6'd40;
			12'd3347 : hue_tab <= 6'd40;
			12'd3348 : hue_tab <= 6'd40;
			12'd3349 : hue_tab <= 6'd40;
			12'd3350 : hue_tab <= 6'd40;
			12'd3351 : hue_tab <= 6'd40;
			12'd3352 : hue_tab <= 6'd40;
			12'd3353 : hue_tab <= 6'd40;
			12'd3354 : hue_tab <= 6'd40;
			12'd3355 : hue_tab <= 6'd40;
			12'd3356 : hue_tab <= 6'd40;
			12'd3357 : hue_tab <= 6'd40;
			12'd3358 : hue_tab <= 6'd40;
			12'd3359 : hue_tab <= 6'd40;
			12'd3360 : hue_tab <= 6'd40;
			12'd3361 : hue_tab <= 6'd40;
			12'd3362 : hue_tab <= 6'd40;
			12'd3363 : hue_tab <= 6'd40;
			12'd3364 : hue_tab <= 6'd40;
			12'd3365 : hue_tab <= 6'd40;
			12'd3366 : hue_tab <= 6'd40;
			12'd3367 : hue_tab <= 6'd40;
			12'd3368 : hue_tab <= 6'd40;
			12'd3369 : hue_tab <= 6'd40;
			12'd3370 : hue_tab <= 6'd40;
			12'd3371 : hue_tab <= 6'd40;
			12'd3372 : hue_tab <= 6'd40;
			12'd3373 : hue_tab <= 6'd40;
			12'd3374 : hue_tab <= 6'd40;
			12'd3375 : hue_tab <= 6'd40;
			12'd3376 : hue_tab <= 6'd40;
			12'd3377 : hue_tab <= 6'd40;
			12'd3378 : hue_tab <= 6'd40;
			12'd3379 : hue_tab <= 6'd40;
			12'd3380 : hue_tab <= 6'd40;
			12'd3381 : hue_tab <= 6'd39;
			12'd3382 : hue_tab <= 6'd38;
			12'd3383 : hue_tab <= 6'd37;
			12'd3384 : hue_tab <= 6'd37;
			12'd3385 : hue_tab <= 6'd36;
			12'd3386 : hue_tab <= 6'd35;
			12'd3387 : hue_tab <= 6'd35;
			12'd3388 : hue_tab <= 6'd34;
			12'd3389 : hue_tab <= 6'd34;
			12'd3390 : hue_tab <= 6'd33;
			12'd3391 : hue_tab <= 6'd33;
			12'd3392 : hue_tab <= 6'd0;
			12'd3393 : hue_tab <= 6'd40;
			12'd3394 : hue_tab <= 6'd40;
			12'd3395 : hue_tab <= 6'd40;
			12'd3396 : hue_tab <= 6'd40;
			12'd3397 : hue_tab <= 6'd40;
			12'd3398 : hue_tab <= 6'd40;
			12'd3399 : hue_tab <= 6'd40;
			12'd3400 : hue_tab <= 6'd40;
			12'd3401 : hue_tab <= 6'd40;
			12'd3402 : hue_tab <= 6'd40;
			12'd3403 : hue_tab <= 6'd40;
			12'd3404 : hue_tab <= 6'd40;
			12'd3405 : hue_tab <= 6'd40;
			12'd3406 : hue_tab <= 6'd40;
			12'd3407 : hue_tab <= 6'd40;
			12'd3408 : hue_tab <= 6'd40;
			12'd3409 : hue_tab <= 6'd40;
			12'd3410 : hue_tab <= 6'd40;
			12'd3411 : hue_tab <= 6'd40;
			12'd3412 : hue_tab <= 6'd40;
			12'd3413 : hue_tab <= 6'd40;
			12'd3414 : hue_tab <= 6'd40;
			12'd3415 : hue_tab <= 6'd40;
			12'd3416 : hue_tab <= 6'd40;
			12'd3417 : hue_tab <= 6'd40;
			12'd3418 : hue_tab <= 6'd40;
			12'd3419 : hue_tab <= 6'd40;
			12'd3420 : hue_tab <= 6'd40;
			12'd3421 : hue_tab <= 6'd40;
			12'd3422 : hue_tab <= 6'd40;
			12'd3423 : hue_tab <= 6'd40;
			12'd3424 : hue_tab <= 6'd40;
			12'd3425 : hue_tab <= 6'd40;
			12'd3426 : hue_tab <= 6'd40;
			12'd3427 : hue_tab <= 6'd40;
			12'd3428 : hue_tab <= 6'd40;
			12'd3429 : hue_tab <= 6'd40;
			12'd3430 : hue_tab <= 6'd40;
			12'd3431 : hue_tab <= 6'd40;
			12'd3432 : hue_tab <= 6'd40;
			12'd3433 : hue_tab <= 6'd40;
			12'd3434 : hue_tab <= 6'd40;
			12'd3435 : hue_tab <= 6'd40;
			12'd3436 : hue_tab <= 6'd40;
			12'd3437 : hue_tab <= 6'd40;
			12'd3438 : hue_tab <= 6'd40;
			12'd3439 : hue_tab <= 6'd40;
			12'd3440 : hue_tab <= 6'd40;
			12'd3441 : hue_tab <= 6'd40;
			12'd3442 : hue_tab <= 6'd40;
			12'd3443 : hue_tab <= 6'd40;
			12'd3444 : hue_tab <= 6'd40;
			12'd3445 : hue_tab <= 6'd40;
			12'd3446 : hue_tab <= 6'd39;
			12'd3447 : hue_tab <= 6'd38;
			12'd3448 : hue_tab <= 6'd37;
			12'd3449 : hue_tab <= 6'd37;
			12'd3450 : hue_tab <= 6'd36;
			12'd3451 : hue_tab <= 6'd35;
			12'd3452 : hue_tab <= 6'd35;
			12'd3453 : hue_tab <= 6'd34;
			12'd3454 : hue_tab <= 6'd34;
			12'd3455 : hue_tab <= 6'd33;
			12'd3456 : hue_tab <= 6'd0;
			12'd3457 : hue_tab <= 6'd40;
			12'd3458 : hue_tab <= 6'd40;
			12'd3459 : hue_tab <= 6'd40;
			12'd3460 : hue_tab <= 6'd40;
			12'd3461 : hue_tab <= 6'd40;
			12'd3462 : hue_tab <= 6'd40;
			12'd3463 : hue_tab <= 6'd40;
			12'd3464 : hue_tab <= 6'd40;
			12'd3465 : hue_tab <= 6'd40;
			12'd3466 : hue_tab <= 6'd40;
			12'd3467 : hue_tab <= 6'd40;
			12'd3468 : hue_tab <= 6'd40;
			12'd3469 : hue_tab <= 6'd40;
			12'd3470 : hue_tab <= 6'd40;
			12'd3471 : hue_tab <= 6'd40;
			12'd3472 : hue_tab <= 6'd40;
			12'd3473 : hue_tab <= 6'd40;
			12'd3474 : hue_tab <= 6'd40;
			12'd3475 : hue_tab <= 6'd40;
			12'd3476 : hue_tab <= 6'd40;
			12'd3477 : hue_tab <= 6'd40;
			12'd3478 : hue_tab <= 6'd40;
			12'd3479 : hue_tab <= 6'd40;
			12'd3480 : hue_tab <= 6'd40;
			12'd3481 : hue_tab <= 6'd40;
			12'd3482 : hue_tab <= 6'd40;
			12'd3483 : hue_tab <= 6'd40;
			12'd3484 : hue_tab <= 6'd40;
			12'd3485 : hue_tab <= 6'd40;
			12'd3486 : hue_tab <= 6'd40;
			12'd3487 : hue_tab <= 6'd40;
			12'd3488 : hue_tab <= 6'd40;
			12'd3489 : hue_tab <= 6'd40;
			12'd3490 : hue_tab <= 6'd40;
			12'd3491 : hue_tab <= 6'd40;
			12'd3492 : hue_tab <= 6'd40;
			12'd3493 : hue_tab <= 6'd40;
			12'd3494 : hue_tab <= 6'd40;
			12'd3495 : hue_tab <= 6'd40;
			12'd3496 : hue_tab <= 6'd40;
			12'd3497 : hue_tab <= 6'd40;
			12'd3498 : hue_tab <= 6'd40;
			12'd3499 : hue_tab <= 6'd40;
			12'd3500 : hue_tab <= 6'd40;
			12'd3501 : hue_tab <= 6'd40;
			12'd3502 : hue_tab <= 6'd40;
			12'd3503 : hue_tab <= 6'd40;
			12'd3504 : hue_tab <= 6'd40;
			12'd3505 : hue_tab <= 6'd40;
			12'd3506 : hue_tab <= 6'd40;
			12'd3507 : hue_tab <= 6'd40;
			12'd3508 : hue_tab <= 6'd40;
			12'd3509 : hue_tab <= 6'd40;
			12'd3510 : hue_tab <= 6'd40;
			12'd3511 : hue_tab <= 6'd39;
			12'd3512 : hue_tab <= 6'd38;
			12'd3513 : hue_tab <= 6'd37;
			12'd3514 : hue_tab <= 6'd37;
			12'd3515 : hue_tab <= 6'd36;
			12'd3516 : hue_tab <= 6'd36;
			12'd3517 : hue_tab <= 6'd35;
			12'd3518 : hue_tab <= 6'd34;
			12'd3519 : hue_tab <= 6'd34;
			12'd3520 : hue_tab <= 6'd0;
			12'd3521 : hue_tab <= 6'd40;
			12'd3522 : hue_tab <= 6'd40;
			12'd3523 : hue_tab <= 6'd40;
			12'd3524 : hue_tab <= 6'd40;
			12'd3525 : hue_tab <= 6'd40;
			12'd3526 : hue_tab <= 6'd40;
			12'd3527 : hue_tab <= 6'd40;
			12'd3528 : hue_tab <= 6'd40;
			12'd3529 : hue_tab <= 6'd40;
			12'd3530 : hue_tab <= 6'd40;
			12'd3531 : hue_tab <= 6'd40;
			12'd3532 : hue_tab <= 6'd40;
			12'd3533 : hue_tab <= 6'd40;
			12'd3534 : hue_tab <= 6'd40;
			12'd3535 : hue_tab <= 6'd40;
			12'd3536 : hue_tab <= 6'd40;
			12'd3537 : hue_tab <= 6'd40;
			12'd3538 : hue_tab <= 6'd40;
			12'd3539 : hue_tab <= 6'd40;
			12'd3540 : hue_tab <= 6'd40;
			12'd3541 : hue_tab <= 6'd40;
			12'd3542 : hue_tab <= 6'd40;
			12'd3543 : hue_tab <= 6'd40;
			12'd3544 : hue_tab <= 6'd40;
			12'd3545 : hue_tab <= 6'd40;
			12'd3546 : hue_tab <= 6'd40;
			12'd3547 : hue_tab <= 6'd40;
			12'd3548 : hue_tab <= 6'd40;
			12'd3549 : hue_tab <= 6'd40;
			12'd3550 : hue_tab <= 6'd40;
			12'd3551 : hue_tab <= 6'd40;
			12'd3552 : hue_tab <= 6'd40;
			12'd3553 : hue_tab <= 6'd40;
			12'd3554 : hue_tab <= 6'd40;
			12'd3555 : hue_tab <= 6'd40;
			12'd3556 : hue_tab <= 6'd40;
			12'd3557 : hue_tab <= 6'd40;
			12'd3558 : hue_tab <= 6'd40;
			12'd3559 : hue_tab <= 6'd40;
			12'd3560 : hue_tab <= 6'd40;
			12'd3561 : hue_tab <= 6'd40;
			12'd3562 : hue_tab <= 6'd40;
			12'd3563 : hue_tab <= 6'd40;
			12'd3564 : hue_tab <= 6'd40;
			12'd3565 : hue_tab <= 6'd40;
			12'd3566 : hue_tab <= 6'd40;
			12'd3567 : hue_tab <= 6'd40;
			12'd3568 : hue_tab <= 6'd40;
			12'd3569 : hue_tab <= 6'd40;
			12'd3570 : hue_tab <= 6'd40;
			12'd3571 : hue_tab <= 6'd40;
			12'd3572 : hue_tab <= 6'd40;
			12'd3573 : hue_tab <= 6'd40;
			12'd3574 : hue_tab <= 6'd40;
			12'd3575 : hue_tab <= 6'd40;
			12'd3576 : hue_tab <= 6'd39;
			12'd3577 : hue_tab <= 6'd38;
			12'd3578 : hue_tab <= 6'd37;
			12'd3579 : hue_tab <= 6'd37;
			12'd3580 : hue_tab <= 6'd36;
			12'd3581 : hue_tab <= 6'd36;
			12'd3582 : hue_tab <= 6'd35;
			12'd3583 : hue_tab <= 6'd34;
			12'd3584 : hue_tab <= 6'd0;
			12'd3585 : hue_tab <= 6'd40;
			12'd3586 : hue_tab <= 6'd40;
			12'd3587 : hue_tab <= 6'd40;
			12'd3588 : hue_tab <= 6'd40;
			12'd3589 : hue_tab <= 6'd40;
			12'd3590 : hue_tab <= 6'd40;
			12'd3591 : hue_tab <= 6'd40;
			12'd3592 : hue_tab <= 6'd40;
			12'd3593 : hue_tab <= 6'd40;
			12'd3594 : hue_tab <= 6'd40;
			12'd3595 : hue_tab <= 6'd40;
			12'd3596 : hue_tab <= 6'd40;
			12'd3597 : hue_tab <= 6'd40;
			12'd3598 : hue_tab <= 6'd40;
			12'd3599 : hue_tab <= 6'd40;
			12'd3600 : hue_tab <= 6'd40;
			12'd3601 : hue_tab <= 6'd40;
			12'd3602 : hue_tab <= 6'd40;
			12'd3603 : hue_tab <= 6'd40;
			12'd3604 : hue_tab <= 6'd40;
			12'd3605 : hue_tab <= 6'd40;
			12'd3606 : hue_tab <= 6'd40;
			12'd3607 : hue_tab <= 6'd40;
			12'd3608 : hue_tab <= 6'd40;
			12'd3609 : hue_tab <= 6'd40;
			12'd3610 : hue_tab <= 6'd40;
			12'd3611 : hue_tab <= 6'd40;
			12'd3612 : hue_tab <= 6'd40;
			12'd3613 : hue_tab <= 6'd40;
			12'd3614 : hue_tab <= 6'd40;
			12'd3615 : hue_tab <= 6'd40;
			12'd3616 : hue_tab <= 6'd40;
			12'd3617 : hue_tab <= 6'd40;
			12'd3618 : hue_tab <= 6'd40;
			12'd3619 : hue_tab <= 6'd40;
			12'd3620 : hue_tab <= 6'd40;
			12'd3621 : hue_tab <= 6'd40;
			12'd3622 : hue_tab <= 6'd40;
			12'd3623 : hue_tab <= 6'd40;
			12'd3624 : hue_tab <= 6'd40;
			12'd3625 : hue_tab <= 6'd40;
			12'd3626 : hue_tab <= 6'd40;
			12'd3627 : hue_tab <= 6'd40;
			12'd3628 : hue_tab <= 6'd40;
			12'd3629 : hue_tab <= 6'd40;
			12'd3630 : hue_tab <= 6'd40;
			12'd3631 : hue_tab <= 6'd40;
			12'd3632 : hue_tab <= 6'd40;
			12'd3633 : hue_tab <= 6'd40;
			12'd3634 : hue_tab <= 6'd40;
			12'd3635 : hue_tab <= 6'd40;
			12'd3636 : hue_tab <= 6'd40;
			12'd3637 : hue_tab <= 6'd40;
			12'd3638 : hue_tab <= 6'd40;
			12'd3639 : hue_tab <= 6'd40;
			12'd3640 : hue_tab <= 6'd40;
			12'd3641 : hue_tab <= 6'd39;
			12'd3642 : hue_tab <= 6'd38;
			12'd3643 : hue_tab <= 6'd37;
			12'd3644 : hue_tab <= 6'd37;
			12'd3645 : hue_tab <= 6'd36;
			12'd3646 : hue_tab <= 6'd36;
			12'd3647 : hue_tab <= 6'd35;
			12'd3648 : hue_tab <= 6'd0;
			12'd3649 : hue_tab <= 6'd40;
			12'd3650 : hue_tab <= 6'd40;
			12'd3651 : hue_tab <= 6'd40;
			12'd3652 : hue_tab <= 6'd40;
			12'd3653 : hue_tab <= 6'd40;
			12'd3654 : hue_tab <= 6'd40;
			12'd3655 : hue_tab <= 6'd40;
			12'd3656 : hue_tab <= 6'd40;
			12'd3657 : hue_tab <= 6'd40;
			12'd3658 : hue_tab <= 6'd40;
			12'd3659 : hue_tab <= 6'd40;
			12'd3660 : hue_tab <= 6'd40;
			12'd3661 : hue_tab <= 6'd40;
			12'd3662 : hue_tab <= 6'd40;
			12'd3663 : hue_tab <= 6'd40;
			12'd3664 : hue_tab <= 6'd40;
			12'd3665 : hue_tab <= 6'd40;
			12'd3666 : hue_tab <= 6'd40;
			12'd3667 : hue_tab <= 6'd40;
			12'd3668 : hue_tab <= 6'd40;
			12'd3669 : hue_tab <= 6'd40;
			12'd3670 : hue_tab <= 6'd40;
			12'd3671 : hue_tab <= 6'd40;
			12'd3672 : hue_tab <= 6'd40;
			12'd3673 : hue_tab <= 6'd40;
			12'd3674 : hue_tab <= 6'd40;
			12'd3675 : hue_tab <= 6'd40;
			12'd3676 : hue_tab <= 6'd40;
			12'd3677 : hue_tab <= 6'd40;
			12'd3678 : hue_tab <= 6'd40;
			12'd3679 : hue_tab <= 6'd40;
			12'd3680 : hue_tab <= 6'd40;
			12'd3681 : hue_tab <= 6'd40;
			12'd3682 : hue_tab <= 6'd40;
			12'd3683 : hue_tab <= 6'd40;
			12'd3684 : hue_tab <= 6'd40;
			12'd3685 : hue_tab <= 6'd40;
			12'd3686 : hue_tab <= 6'd40;
			12'd3687 : hue_tab <= 6'd40;
			12'd3688 : hue_tab <= 6'd40;
			12'd3689 : hue_tab <= 6'd40;
			12'd3690 : hue_tab <= 6'd40;
			12'd3691 : hue_tab <= 6'd40;
			12'd3692 : hue_tab <= 6'd40;
			12'd3693 : hue_tab <= 6'd40;
			12'd3694 : hue_tab <= 6'd40;
			12'd3695 : hue_tab <= 6'd40;
			12'd3696 : hue_tab <= 6'd40;
			12'd3697 : hue_tab <= 6'd40;
			12'd3698 : hue_tab <= 6'd40;
			12'd3699 : hue_tab <= 6'd40;
			12'd3700 : hue_tab <= 6'd40;
			12'd3701 : hue_tab <= 6'd40;
			12'd3702 : hue_tab <= 6'd40;
			12'd3703 : hue_tab <= 6'd40;
			12'd3704 : hue_tab <= 6'd40;
			12'd3705 : hue_tab <= 6'd40;
			12'd3706 : hue_tab <= 6'd39;
			12'd3707 : hue_tab <= 6'd38;
			12'd3708 : hue_tab <= 6'd38;
			12'd3709 : hue_tab <= 6'd37;
			12'd3710 : hue_tab <= 6'd36;
			12'd3711 : hue_tab <= 6'd36;
			12'd3712 : hue_tab <= 6'd0;
			12'd3713 : hue_tab <= 6'd40;
			12'd3714 : hue_tab <= 6'd40;
			12'd3715 : hue_tab <= 6'd40;
			12'd3716 : hue_tab <= 6'd40;
			12'd3717 : hue_tab <= 6'd40;
			12'd3718 : hue_tab <= 6'd40;
			12'd3719 : hue_tab <= 6'd40;
			12'd3720 : hue_tab <= 6'd40;
			12'd3721 : hue_tab <= 6'd40;
			12'd3722 : hue_tab <= 6'd40;
			12'd3723 : hue_tab <= 6'd40;
			12'd3724 : hue_tab <= 6'd40;
			12'd3725 : hue_tab <= 6'd40;
			12'd3726 : hue_tab <= 6'd40;
			12'd3727 : hue_tab <= 6'd40;
			12'd3728 : hue_tab <= 6'd40;
			12'd3729 : hue_tab <= 6'd40;
			12'd3730 : hue_tab <= 6'd40;
			12'd3731 : hue_tab <= 6'd40;
			12'd3732 : hue_tab <= 6'd40;
			12'd3733 : hue_tab <= 6'd40;
			12'd3734 : hue_tab <= 6'd40;
			12'd3735 : hue_tab <= 6'd40;
			12'd3736 : hue_tab <= 6'd40;
			12'd3737 : hue_tab <= 6'd40;
			12'd3738 : hue_tab <= 6'd40;
			12'd3739 : hue_tab <= 6'd40;
			12'd3740 : hue_tab <= 6'd40;
			12'd3741 : hue_tab <= 6'd40;
			12'd3742 : hue_tab <= 6'd40;
			12'd3743 : hue_tab <= 6'd40;
			12'd3744 : hue_tab <= 6'd40;
			12'd3745 : hue_tab <= 6'd40;
			12'd3746 : hue_tab <= 6'd40;
			12'd3747 : hue_tab <= 6'd40;
			12'd3748 : hue_tab <= 6'd40;
			12'd3749 : hue_tab <= 6'd40;
			12'd3750 : hue_tab <= 6'd40;
			12'd3751 : hue_tab <= 6'd40;
			12'd3752 : hue_tab <= 6'd40;
			12'd3753 : hue_tab <= 6'd40;
			12'd3754 : hue_tab <= 6'd40;
			12'd3755 : hue_tab <= 6'd40;
			12'd3756 : hue_tab <= 6'd40;
			12'd3757 : hue_tab <= 6'd40;
			12'd3758 : hue_tab <= 6'd40;
			12'd3759 : hue_tab <= 6'd40;
			12'd3760 : hue_tab <= 6'd40;
			12'd3761 : hue_tab <= 6'd40;
			12'd3762 : hue_tab <= 6'd40;
			12'd3763 : hue_tab <= 6'd40;
			12'd3764 : hue_tab <= 6'd40;
			12'd3765 : hue_tab <= 6'd40;
			12'd3766 : hue_tab <= 6'd40;
			12'd3767 : hue_tab <= 6'd40;
			12'd3768 : hue_tab <= 6'd40;
			12'd3769 : hue_tab <= 6'd40;
			12'd3770 : hue_tab <= 6'd40;
			12'd3771 : hue_tab <= 6'd39;
			12'd3772 : hue_tab <= 6'd38;
			12'd3773 : hue_tab <= 6'd38;
			12'd3774 : hue_tab <= 6'd37;
			12'd3775 : hue_tab <= 6'd36;
			12'd3776 : hue_tab <= 6'd0;
			12'd3777 : hue_tab <= 6'd40;
			12'd3778 : hue_tab <= 6'd40;
			12'd3779 : hue_tab <= 6'd40;
			12'd3780 : hue_tab <= 6'd40;
			12'd3781 : hue_tab <= 6'd40;
			12'd3782 : hue_tab <= 6'd40;
			12'd3783 : hue_tab <= 6'd40;
			12'd3784 : hue_tab <= 6'd40;
			12'd3785 : hue_tab <= 6'd40;
			12'd3786 : hue_tab <= 6'd40;
			12'd3787 : hue_tab <= 6'd40;
			12'd3788 : hue_tab <= 6'd40;
			12'd3789 : hue_tab <= 6'd40;
			12'd3790 : hue_tab <= 6'd40;
			12'd3791 : hue_tab <= 6'd40;
			12'd3792 : hue_tab <= 6'd40;
			12'd3793 : hue_tab <= 6'd40;
			12'd3794 : hue_tab <= 6'd40;
			12'd3795 : hue_tab <= 6'd40;
			12'd3796 : hue_tab <= 6'd40;
			12'd3797 : hue_tab <= 6'd40;
			12'd3798 : hue_tab <= 6'd40;
			12'd3799 : hue_tab <= 6'd40;
			12'd3800 : hue_tab <= 6'd40;
			12'd3801 : hue_tab <= 6'd40;
			12'd3802 : hue_tab <= 6'd40;
			12'd3803 : hue_tab <= 6'd40;
			12'd3804 : hue_tab <= 6'd40;
			12'd3805 : hue_tab <= 6'd40;
			12'd3806 : hue_tab <= 6'd40;
			12'd3807 : hue_tab <= 6'd40;
			12'd3808 : hue_tab <= 6'd40;
			12'd3809 : hue_tab <= 6'd40;
			12'd3810 : hue_tab <= 6'd40;
			12'd3811 : hue_tab <= 6'd40;
			12'd3812 : hue_tab <= 6'd40;
			12'd3813 : hue_tab <= 6'd40;
			12'd3814 : hue_tab <= 6'd40;
			12'd3815 : hue_tab <= 6'd40;
			12'd3816 : hue_tab <= 6'd40;
			12'd3817 : hue_tab <= 6'd40;
			12'd3818 : hue_tab <= 6'd40;
			12'd3819 : hue_tab <= 6'd40;
			12'd3820 : hue_tab <= 6'd40;
			12'd3821 : hue_tab <= 6'd40;
			12'd3822 : hue_tab <= 6'd40;
			12'd3823 : hue_tab <= 6'd40;
			12'd3824 : hue_tab <= 6'd40;
			12'd3825 : hue_tab <= 6'd40;
			12'd3826 : hue_tab <= 6'd40;
			12'd3827 : hue_tab <= 6'd40;
			12'd3828 : hue_tab <= 6'd40;
			12'd3829 : hue_tab <= 6'd40;
			12'd3830 : hue_tab <= 6'd40;
			12'd3831 : hue_tab <= 6'd40;
			12'd3832 : hue_tab <= 6'd40;
			12'd3833 : hue_tab <= 6'd40;
			12'd3834 : hue_tab <= 6'd40;
			12'd3835 : hue_tab <= 6'd40;
			12'd3836 : hue_tab <= 6'd39;
			12'd3837 : hue_tab <= 6'd38;
			12'd3838 : hue_tab <= 6'd38;
			12'd3839 : hue_tab <= 6'd37;
			12'd3840 : hue_tab <= 6'd0;
			12'd3841 : hue_tab <= 6'd40;
			12'd3842 : hue_tab <= 6'd40;
			12'd3843 : hue_tab <= 6'd40;
			12'd3844 : hue_tab <= 6'd40;
			12'd3845 : hue_tab <= 6'd40;
			12'd3846 : hue_tab <= 6'd40;
			12'd3847 : hue_tab <= 6'd40;
			12'd3848 : hue_tab <= 6'd40;
			12'd3849 : hue_tab <= 6'd40;
			12'd3850 : hue_tab <= 6'd40;
			12'd3851 : hue_tab <= 6'd40;
			12'd3852 : hue_tab <= 6'd40;
			12'd3853 : hue_tab <= 6'd40;
			12'd3854 : hue_tab <= 6'd40;
			12'd3855 : hue_tab <= 6'd40;
			12'd3856 : hue_tab <= 6'd40;
			12'd3857 : hue_tab <= 6'd40;
			12'd3858 : hue_tab <= 6'd40;
			12'd3859 : hue_tab <= 6'd40;
			12'd3860 : hue_tab <= 6'd40;
			12'd3861 : hue_tab <= 6'd40;
			12'd3862 : hue_tab <= 6'd40;
			12'd3863 : hue_tab <= 6'd40;
			12'd3864 : hue_tab <= 6'd40;
			12'd3865 : hue_tab <= 6'd40;
			12'd3866 : hue_tab <= 6'd40;
			12'd3867 : hue_tab <= 6'd40;
			12'd3868 : hue_tab <= 6'd40;
			12'd3869 : hue_tab <= 6'd40;
			12'd3870 : hue_tab <= 6'd40;
			12'd3871 : hue_tab <= 6'd40;
			12'd3872 : hue_tab <= 6'd40;
			12'd3873 : hue_tab <= 6'd40;
			12'd3874 : hue_tab <= 6'd40;
			12'd3875 : hue_tab <= 6'd40;
			12'd3876 : hue_tab <= 6'd40;
			12'd3877 : hue_tab <= 6'd40;
			12'd3878 : hue_tab <= 6'd40;
			12'd3879 : hue_tab <= 6'd40;
			12'd3880 : hue_tab <= 6'd40;
			12'd3881 : hue_tab <= 6'd40;
			12'd3882 : hue_tab <= 6'd40;
			12'd3883 : hue_tab <= 6'd40;
			12'd3884 : hue_tab <= 6'd40;
			12'd3885 : hue_tab <= 6'd40;
			12'd3886 : hue_tab <= 6'd40;
			12'd3887 : hue_tab <= 6'd40;
			12'd3888 : hue_tab <= 6'd40;
			12'd3889 : hue_tab <= 6'd40;
			12'd3890 : hue_tab <= 6'd40;
			12'd3891 : hue_tab <= 6'd40;
			12'd3892 : hue_tab <= 6'd40;
			12'd3893 : hue_tab <= 6'd40;
			12'd3894 : hue_tab <= 6'd40;
			12'd3895 : hue_tab <= 6'd40;
			12'd3896 : hue_tab <= 6'd40;
			12'd3897 : hue_tab <= 6'd40;
			12'd3898 : hue_tab <= 6'd40;
			12'd3899 : hue_tab <= 6'd40;
			12'd3900 : hue_tab <= 6'd40;
			12'd3901 : hue_tab <= 6'd39;
			12'd3902 : hue_tab <= 6'd38;
			12'd3903 : hue_tab <= 6'd38;
			12'd3904 : hue_tab <= 6'd0;
			12'd3905 : hue_tab <= 6'd40;
			12'd3906 : hue_tab <= 6'd40;
			12'd3907 : hue_tab <= 6'd40;
			12'd3908 : hue_tab <= 6'd40;
			12'd3909 : hue_tab <= 6'd40;
			12'd3910 : hue_tab <= 6'd40;
			12'd3911 : hue_tab <= 6'd40;
			12'd3912 : hue_tab <= 6'd40;
			12'd3913 : hue_tab <= 6'd40;
			12'd3914 : hue_tab <= 6'd40;
			12'd3915 : hue_tab <= 6'd40;
			12'd3916 : hue_tab <= 6'd40;
			12'd3917 : hue_tab <= 6'd40;
			12'd3918 : hue_tab <= 6'd40;
			12'd3919 : hue_tab <= 6'd40;
			12'd3920 : hue_tab <= 6'd40;
			12'd3921 : hue_tab <= 6'd40;
			12'd3922 : hue_tab <= 6'd40;
			12'd3923 : hue_tab <= 6'd40;
			12'd3924 : hue_tab <= 6'd40;
			12'd3925 : hue_tab <= 6'd40;
			12'd3926 : hue_tab <= 6'd40;
			12'd3927 : hue_tab <= 6'd40;
			12'd3928 : hue_tab <= 6'd40;
			12'd3929 : hue_tab <= 6'd40;
			12'd3930 : hue_tab <= 6'd40;
			12'd3931 : hue_tab <= 6'd40;
			12'd3932 : hue_tab <= 6'd40;
			12'd3933 : hue_tab <= 6'd40;
			12'd3934 : hue_tab <= 6'd40;
			12'd3935 : hue_tab <= 6'd40;
			12'd3936 : hue_tab <= 6'd40;
			12'd3937 : hue_tab <= 6'd40;
			12'd3938 : hue_tab <= 6'd40;
			12'd3939 : hue_tab <= 6'd40;
			12'd3940 : hue_tab <= 6'd40;
			12'd3941 : hue_tab <= 6'd40;
			12'd3942 : hue_tab <= 6'd40;
			12'd3943 : hue_tab <= 6'd40;
			12'd3944 : hue_tab <= 6'd40;
			12'd3945 : hue_tab <= 6'd40;
			12'd3946 : hue_tab <= 6'd40;
			12'd3947 : hue_tab <= 6'd40;
			12'd3948 : hue_tab <= 6'd40;
			12'd3949 : hue_tab <= 6'd40;
			12'd3950 : hue_tab <= 6'd40;
			12'd3951 : hue_tab <= 6'd40;
			12'd3952 : hue_tab <= 6'd40;
			12'd3953 : hue_tab <= 6'd40;
			12'd3954 : hue_tab <= 6'd40;
			12'd3955 : hue_tab <= 6'd40;
			12'd3956 : hue_tab <= 6'd40;
			12'd3957 : hue_tab <= 6'd40;
			12'd3958 : hue_tab <= 6'd40;
			12'd3959 : hue_tab <= 6'd40;
			12'd3960 : hue_tab <= 6'd40;
			12'd3961 : hue_tab <= 6'd40;
			12'd3962 : hue_tab <= 6'd40;
			12'd3963 : hue_tab <= 6'd40;
			12'd3964 : hue_tab <= 6'd40;
			12'd3965 : hue_tab <= 6'd40;
			12'd3966 : hue_tab <= 6'd39;
			12'd3967 : hue_tab <= 6'd38;
			12'd3968 : hue_tab <= 6'd0;
			12'd3969 : hue_tab <= 6'd40;
			12'd3970 : hue_tab <= 6'd40;
			12'd3971 : hue_tab <= 6'd40;
			12'd3972 : hue_tab <= 6'd40;
			12'd3973 : hue_tab <= 6'd40;
			12'd3974 : hue_tab <= 6'd40;
			12'd3975 : hue_tab <= 6'd40;
			12'd3976 : hue_tab <= 6'd40;
			12'd3977 : hue_tab <= 6'd40;
			12'd3978 : hue_tab <= 6'd40;
			12'd3979 : hue_tab <= 6'd40;
			12'd3980 : hue_tab <= 6'd40;
			12'd3981 : hue_tab <= 6'd40;
			12'd3982 : hue_tab <= 6'd40;
			12'd3983 : hue_tab <= 6'd40;
			12'd3984 : hue_tab <= 6'd40;
			12'd3985 : hue_tab <= 6'd40;
			12'd3986 : hue_tab <= 6'd40;
			12'd3987 : hue_tab <= 6'd40;
			12'd3988 : hue_tab <= 6'd40;
			12'd3989 : hue_tab <= 6'd40;
			12'd3990 : hue_tab <= 6'd40;
			12'd3991 : hue_tab <= 6'd40;
			12'd3992 : hue_tab <= 6'd40;
			12'd3993 : hue_tab <= 6'd40;
			12'd3994 : hue_tab <= 6'd40;
			12'd3995 : hue_tab <= 6'd40;
			12'd3996 : hue_tab <= 6'd40;
			12'd3997 : hue_tab <= 6'd40;
			12'd3998 : hue_tab <= 6'd40;
			12'd3999 : hue_tab <= 6'd40;
			12'd4000 : hue_tab <= 6'd40;
			12'd4001 : hue_tab <= 6'd40;
			12'd4002 : hue_tab <= 6'd40;
			12'd4003 : hue_tab <= 6'd40;
			12'd4004 : hue_tab <= 6'd40;
			12'd4005 : hue_tab <= 6'd40;
			12'd4006 : hue_tab <= 6'd40;
			12'd4007 : hue_tab <= 6'd40;
			12'd4008 : hue_tab <= 6'd40;
			12'd4009 : hue_tab <= 6'd40;
			12'd4010 : hue_tab <= 6'd40;
			12'd4011 : hue_tab <= 6'd40;
			12'd4012 : hue_tab <= 6'd40;
			12'd4013 : hue_tab <= 6'd40;
			12'd4014 : hue_tab <= 6'd40;
			12'd4015 : hue_tab <= 6'd40;
			12'd4016 : hue_tab <= 6'd40;
			12'd4017 : hue_tab <= 6'd40;
			12'd4018 : hue_tab <= 6'd40;
			12'd4019 : hue_tab <= 6'd40;
			12'd4020 : hue_tab <= 6'd40;
			12'd4021 : hue_tab <= 6'd40;
			12'd4022 : hue_tab <= 6'd40;
			12'd4023 : hue_tab <= 6'd40;
			12'd4024 : hue_tab <= 6'd40;
			12'd4025 : hue_tab <= 6'd40;
			12'd4026 : hue_tab <= 6'd40;
			12'd4027 : hue_tab <= 6'd40;
			12'd4028 : hue_tab <= 6'd40;
			12'd4029 : hue_tab <= 6'd40;
			12'd4030 : hue_tab <= 6'd40;
			12'd4031 : hue_tab <= 6'd39;
			12'd4032 : hue_tab <= 6'd0;
			12'd4033 : hue_tab <= 6'd40;
			12'd4034 : hue_tab <= 6'd40;
			12'd4035 : hue_tab <= 6'd40;
			12'd4036 : hue_tab <= 6'd40;
			12'd4037 : hue_tab <= 6'd40;
			12'd4038 : hue_tab <= 6'd40;
			12'd4039 : hue_tab <= 6'd40;
			12'd4040 : hue_tab <= 6'd40;
			12'd4041 : hue_tab <= 6'd40;
			12'd4042 : hue_tab <= 6'd40;
			12'd4043 : hue_tab <= 6'd40;
			12'd4044 : hue_tab <= 6'd40;
			12'd4045 : hue_tab <= 6'd40;
			12'd4046 : hue_tab <= 6'd40;
			12'd4047 : hue_tab <= 6'd40;
			12'd4048 : hue_tab <= 6'd40;
			12'd4049 : hue_tab <= 6'd40;
			12'd4050 : hue_tab <= 6'd40;
			12'd4051 : hue_tab <= 6'd40;
			12'd4052 : hue_tab <= 6'd40;
			12'd4053 : hue_tab <= 6'd40;
			12'd4054 : hue_tab <= 6'd40;
			12'd4055 : hue_tab <= 6'd40;
			12'd4056 : hue_tab <= 6'd40;
			12'd4057 : hue_tab <= 6'd40;
			12'd4058 : hue_tab <= 6'd40;
			12'd4059 : hue_tab <= 6'd40;
			12'd4060 : hue_tab <= 6'd40;
			12'd4061 : hue_tab <= 6'd40;
			12'd4062 : hue_tab <= 6'd40;
			12'd4063 : hue_tab <= 6'd40;
			12'd4064 : hue_tab <= 6'd40;
			12'd4065 : hue_tab <= 6'd40;
			12'd4066 : hue_tab <= 6'd40;
			12'd4067 : hue_tab <= 6'd40;
			12'd4068 : hue_tab <= 6'd40;
			12'd4069 : hue_tab <= 6'd40;
			12'd4070 : hue_tab <= 6'd40;
			12'd4071 : hue_tab <= 6'd40;
			12'd4072 : hue_tab <= 6'd40;
			12'd4073 : hue_tab <= 6'd40;
			12'd4074 : hue_tab <= 6'd40;
			12'd4075 : hue_tab <= 6'd40;
			12'd4076 : hue_tab <= 6'd40;
			12'd4077 : hue_tab <= 6'd40;
			12'd4078 : hue_tab <= 6'd40;
			12'd4079 : hue_tab <= 6'd40;
			12'd4080 : hue_tab <= 6'd40;
			12'd4081 : hue_tab <= 6'd40;
			12'd4082 : hue_tab <= 6'd40;
			12'd4083 : hue_tab <= 6'd40;
			12'd4084 : hue_tab <= 6'd40;
			12'd4085 : hue_tab <= 6'd40;
			12'd4086 : hue_tab <= 6'd40;
			12'd4087 : hue_tab <= 6'd40;
			12'd4088 : hue_tab <= 6'd40;
			12'd4089 : hue_tab <= 6'd40;
			12'd4090 : hue_tab <= 6'd40;
			12'd4091 : hue_tab <= 6'd40;
			12'd4092 : hue_tab <= 6'd40;
			12'd4093 : hue_tab <= 6'd40;
			12'd4094 : hue_tab <= 6'd40;
			12'd4095 : hue_tab <= 6'd40;
	endcase
end

reg [3:0] last_hue_ofs, last2_hue_ofs;
reg last_sub, last2_sub;
always @(posedge clk) begin
	last_hue_ofs <= hue_ofs;
	last2_hue_ofs <= last_hue_ofs;
	last_sub <= sub;
	last2_sub <= last_sub;
	hue <= {last2_hue_ofs,4'h0} + (last2_sub ? -hue_tab : hue_tab);
end

endmodule