module int_test(address, instruction, clk);
input [7:0] address;
output [15:0] instruction;
input clk;
RAMB4_S16 ram_256_x_16(
	.DI  (16'b0),
	.EN (1'b1),
	.WE (1'b0),
	.RST (1'b0),
	.CLK (clk),
	.ADDR(address),
	.DO (instruction)
);
// synthesis translate_off
defparam ram_256_x_16.INIT_00 = 256'h0000000000000000000000000000810332FF950560010007E202803002AA0A00;
defparam ram_256_x_16.INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_256_x_16.INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_256_x_16.INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_256_x_16.INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_256_x_16.INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_256_x_16.INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_256_x_16.INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_256_x_16.INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_256_x_16.INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_256_x_16.INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_256_x_16.INIT_0B = 256'h000000000000000000000000000000000000000000000000000080F0EA044A01;
defparam ram_256_x_16.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_256_x_16.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_256_x_16.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ram_256_x_16.INIT_0F = 256'h81B0000000000000000000000000000000000000000000000000000000000000;
// synthesis translate_on
// synthesis attribute INIT_00 of ram_256_x_16 is "0000000000000000000000000000810332FF950560010007E202803002AA0A00"
// synthesis attribute INIT_01 of ram_256_x_16 is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_02 of ram_256_x_16 is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_03 of ram_256_x_16 is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_04 of ram_256_x_16 is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_05 of ram_256_x_16 is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_06 of ram_256_x_16 is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_07 of ram_256_x_16 is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_08 of ram_256_x_16 is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_09 of ram_256_x_16 is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_0A of ram_256_x_16 is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_0B of ram_256_x_16 is "000000000000000000000000000000000000000000000000000080F0EA044A01"
// synthesis attribute INIT_0C of ram_256_x_16 is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_0D of ram_256_x_16 is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_0E of ram_256_x_16 is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_0F of ram_256_x_16 is "81B0000000000000000000000000000000000000000000000000000000000000"
endmodule
