`define WIDTH 5